BZh91AY&SY��w> m_�Px����߰����P^9lwɐD@�B��F�����SG�SA� =&����̦�	�4�14dd���d�S"��MM�M 4  40`��`ѐ��&��D��h��=(�����#LOP�I$���
�"hI���	>�������}�{)��XBjT_FN;�1"�m�CH���t�o>�t\�\��&[S!emƫmI�����&a�-Ͷr�'h��Q"6��O��g�$B�1�i��A�v�E	�1n�]�ÿ��M�fM��{m�r�����k����~b�X<IP�.;P���c��ad�=�L"֘��E@�6�N��Wpp���̦��r%�j��N���_)�ns�X�l(��XK&V/�2c��E�v�w������P��P5y�H�W�b\���Xk$N.M�t"���Ү�s����������$�HAd����LG�w�h�Zwۺ%M��|6���2DP�%H����J�SE�չ �G}�Yޜ�&L.�:ַ���,��4=}����@�~�w��ЈD[�<�����C#3��  �T��3�XJvO̢!x`����O�����*�@��RN{��H<i((z�~�Y��(�3�++���o�r����f��@�廬MI��ڬ��%
W���^�t��	jӖ��1�:�=����fb�F�SQ^�Úi��K���FI�����q�D�5Z�9ƹt�w�tfl��W㮂=T��@J%B���zTD��V�M)��e�Z��|��jT����^-��5b_�4.>��2�8R$��bWFX�*.��%8�dG�">�۳b`�ޜǅjE��R�Аnw��=,tю����Y!�b��.��V�W&(!IE�61��}���"XvuS�f�Y���4��<�x�9N'��r�L1@:"�4Zɢ���=m����Nıi �5/�ْ0J��� ��G���՜QZ$�����3��y��
7i\.	���QBQ
��7f�`9�E�����O��'����9��0���������{!5��B5���!��	�MҾS�w6�A��.�iX�����%^@ld��9�fN�0���de=T�=�e�}t���tTX�	aZ�V]3�p��S���X1
�I͏n4f�R��̪�<��qm�v�tb<&���D��m`rT���!Z���A}Y�jS(�0��8< ����2)&b?\V����$Zɒ.��5���w$S�	
��s�