BZh91AY&SYV�B t߀Px����߰����`-��Np*T����	�Bz5Oh��Sh��~�S�zh��z�T��)        `LM&L�LM21001E =@��� d  4 ���a2dɑ��4�# C �"��F�?T�6�E=1@���&��	���L`���T�Q(Y�=��D>��xe@O�D#P1=нP{�	�$N��q������ؤ���d}�@I�.�����8��9|��JL����2��-9)�0�L��l��΃��C燩��oX��EFr�!���N.'��6&� `^�WAq�7Q��}9f�!2`oL���{?cיw�/��KM�ps�����DV�	fR2z��U#[l+��`�g����2.h�A��Н�k�a��e���!�&�'!����3zD��/���oE̲��Bg��E{�D'��X���+|��;��^ؙ�d8�:5d21-1�L-��� a��H�ނfJ�0�A
��;�A�����)ÑL3��C�D�JX��@
��HAIi��Sy$<e�Q�$�
�L�Zf������w8�6�ER�7�N��Q�"�-J�0B��BL�T%�Af�F	k+,@����f�҅[9v��S{��s�ϯ���ĐH$�	$� v�o��#ϳmE�ԬC#��`��X|���*�Z�-DR�`7��u���J��B/t�(헙l�T�ex_��!3 U��ƿ�����NUUՆ{��˄����<|`_g�����k���4�������j�SHA�v���ҫ��@�R[L
<h#×��#ƍeoYU�t���Y��`�iZ6]�8Ϳ����0��̐���`��;��7�7")G�P���o�4zԨ�n]{W�cT�y�� ��/&1�h�X�=��x����k.D-O6o��]���v�t�O}!d�w�''�|"���G^Ǆ0�S �- ̊Q\ �F_V8�E��bi�j=�p��B[��v�uv^^�6����"�l�ER�P__rB
H�����s��.FY��R���4��s���ry���Y���]8i�Vi!��`��`�@|ij���bB�C�{�i���G>��h�>�2�\��sA�Q�������I�uhy�Z��8�2*!�Xr�rܤa�]��� �m��aa.0sl�xR�`���L�QtĖhL���� D ��v�t�6���:Bm�$�����W������s7|�Y�ͮ�|�`�Sd�#��t�}��Bo��D�aiC��a7��.z=����Bz����^�a�j��b	8vZ+!vQ5�vF0�4�&�f3������T���gb��4�HLyA�6�	&�#]��s;
�QsO��ѠP��������:sI���E���U�o�@�ö�r�Ģ�%7#�8�x\4�=�����˾�*���ѥvr_��H�

��C�