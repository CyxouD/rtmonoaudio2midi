BZh91AY&SY�+r' p_�Px����߰����`_,�q�@�UQ	$I�4��O&jl��aOQ��Pi���z��SR�       4d���`F�b0L�`��B ����@   @sFLL LFi�#ɀF		�b	���F��Tɉ�F����� C�t�V$L%I���x�HA����Se�Q!P������4	V6���*��wo\=Zp�!%��L)����	߾N�Jm�[�!��;�M��;@2e��!Qޒ�96�C�����_W=5��:t���i[k)�����f8���� �(��$���$	)��!�����$�������,�n���}�qZ�6{��GC�EϠ�v��	���
6A��.�_v��U�J<� D�&�B� ���\+l8mhm]O5���gNj���(��1����jd�YdX���<�K�:���O3&��^v����]f0�AA�J�;�@�3bmRĒ!ڥQ(�̻iNb�V&nL,�Y�L,*�
�-v��a@���M��o$��+�B���Ur^>F�fH�2��a�3BBf[�r�&j�)g���o���ȼ����ZPϨd��	2�1)R&E�+l)R���"vM�e�ۏ��g �� L �{���d��uy���%㈫$��P*Y6i}g�c����性����X�\������p]�+�\�Y�zC��f9������Q�J5U����޶����gd��>O�_�.�*�_'���q+�OJ�B7��xx_�	��+�O7����M�-�{N���V2l��b׿.A�������Ɔ�x��˟h��Swۭc���S�9��m6A�Q�3z�f��E��.���:q̚��L7�"��$���3BD�m��s8�VBV���n�R�cm�L��^[�%F��y�g�p>���H�� �&���:ZF�| �p��G���Ƞ�RI"X�ݥ3M��cJ�Pd1�ÎؒoI�\t`�T^�B
j�:�܈�ӯj`� ����Q$]�2�l�Q�@��̐-��)2l־E��=�êd�Zn��L��B
h���=R{Ϸ0>�+�>:an�u�Mf��k�Ԑ���\@���xW���`>�tE�4�E�URz���i�4�%�"Խ�fHD�e)' �|#}/���(�t�����3c�r*A
�y.�{�r(�i2� Ϩ�vb/��h�׃ǳ�S�^�y��hoTC��ˬl<�g�6�G�y_bV�B�zi����@a�!��|�殣vN�`�����\����Gn�zOn�t`���<Ҭ�FV�$���EuQ� �Q��|�$ �� �R�9�Y�6B��eVy�᫞��-bAp��+�$n��d��ֽ͓�8AןI\��Ў}GOL�`�b6�&Uz,K�+�is�32d�k���ܑN$$
܉�