BZh91AY&SYiHG _�Px����߰����P��n�▌�j�$����i3@��4&'��yF����h5OȘ�J�       �	4B��hz�#���h4 ɵ�& �4d40	�10�@ !I���OdО�S��=P0 �	�$��I HK�@��>K`���`��`�#�50�$+��G&iaf�=KW��@G�+�MIc�8
t��ޔ;5��y]k%���i��;��4�3Mh��NYA#�9����ΙrA�(��*���\���>�QL��M��W]�z���j!���~�ۤ\�)�!��(c��u��gF/".0Y�0��`��J�i����e�� v'm
� T��#���Id���wA3o���5��0"�7L����E������P����)I�qm �-I9�/�Y"t��cI��4��: ��20C�l�l���8�;ݻc6͇����b���U?�.�>C[llm��m� �p�ԧ���=�k+է��%���v+�c2i�T6Z9�#����-,�Z&(1w���)@�PW0���O�4�c5�5���6��R�ǆ��aܹ�{�,��o�W������~��/��w�ɰrKB�������J��Ĥ<��	��M�O�ɇ�5%/Y��j9۾%l��jÞ���U�C� �!X846?����'�������N��˘�c�=|Y4�A�y�q�nk3T4
�:~���	�'�m��R��,v_Ʒs�J�P�Ƶ�nX�Y�u���m@�t���P4wZR�h�h ܖ��N����	p�@s����d�" !��~i��W��j�1���Sz�c��k��^O�o��={��# �"�)Y�S^��1��C�)�b��-x��H���c(�m�s@}K���Sk�c�9��aϽ��4��ƊSY����B�>+�8#�}w��{� �|� �j�HV�ꪓ���tHfI;��
����$E ��N����2*��Y^%AN
%�]�	�����r�'��"h�6���J����f)o�3���4�TN=��=,�9�u�z`�+Y#�l5�R�X�C�Rؙu��{@D�h�͞E*�w���%nF�9$���Ió⬄�H �?|%�u�Y�-���Z���$n�2U\%�`��C}ٺ �0<M�c�r��
5 d9Y煮[.��!k
� �I"��m���S����l,]�g �^Rz�
.F<\��@��do1��b?|7=���$\ɒ3��v���H�
�)�