BZh91AY&SY�@d� J_�Px����߰����`/��u�U$����ҟ��c<�2����C M���T��IH L �4� ���#ja d�0�@�Ms F	�0M`�Ls F	�0M`�L$D �h���́&��M���Fj ɴD�S�zI�$E$	:BD�8�w�����ʌ��`�����GƂB1"�m�!�U��ut�_X�ҷ�,� ����k��Ts̬��e�T�K��l��l�d٪3e�Ɏ>n8�#1PhY�*���؃HY˔����	h���?����$� f?t�A���Ǘ���+@�H��qv��CG[�\5%�p��q�"D���n���,btרa(���р�;d;�&��oƐ�Aڅ;R��D���;�A-H�i,tS�&s���]5i��! ei6ҐDj��� j��v,�l�F<ja���Zm
w��C�����*4�epe;x���jo���Me�6f	ɚj}�chd�Fa���J�Ijm�A#0�!ӵ�65�J3�d��;�	�.Z��8Ͱc���1új�}W� �3r��)��]���~/�v�cco��m�hA۷�O������Y��Y�θ���a��i1��xDL2���<XbҖ�m�L\�s
���]�/j����1$�B����P���=}2��9�8H��?"����������/|�WQ�V;�� �g����c��0�$Ӆ	�g&ۣ��bMQT����w�J��㗠Aȭ����;� ��_p�v��A��`7������.Lh�Rާ�H��i�B8�כJ�˂�� ���]L~/�i�l��a��>�u$D�,�]yߧ�JQOˊ�!%�YJ�y	Qa2t4�����@�CD0�$Z��-)�k|��*��p;hGQ��i*VH�[�Rf���5��cv��Ħ���eE��{� ��H����A2��nT[UpE��O�ۂa����J	d��-�-����W���b��ܴ'%��-u�� A]�Ǯ^�����N�5���nШ����i!� ��`�8щ�{��(��Qqz�
�����1��#2�؜�S�]�"(*^�8~p�Z�`+��*��PE	��f�r� �P�ݷ|}9��9}�6]�csƭ���*��#O��PAS5��u��`�[G�'��د���GJd��-A`5� u>�!A�����,ɞjU�T�UͨT��]��E�'��ᦺ��^�G��/��n��2'v9��z���E��jv��;a�����A�t,��E�͸b���D��4�H��ؗ�ĵk"[U,�4�ǁF5%���a��@����e5K�m�f9��/d��>�����)��&