BZh91AY&SY �� �߀Px����߰����P��m���lFf�ВAh#*��)榨�OSʛQ�SڍFG��yC����4�T4 22bddbh20�H��L���1��@�� mOP2dɈ��	�����$Q1b���G�➚�<���   �$eם$�1"� HK�@��:�l���Q�`�#hjG��bꠐ�"lmA�M�msv��m�6El٤�~`���������E�f��BH)߉s1ʒ�&).!Ù�oP�2�m��Ҥ���X�k���;̌	h.���./	���!BX�HEb�0Ύ=Ǐ\� �``���=z���ڻ��wy�A����Kp�/�R�U�����/�𴨐�:
� lM�*E&k��݈H��;�bɥ���$$!��!����RB��\jQ*�)p��J����qW[]
d ���o�Y[�E�R�(V���E=]�(UP���!�CC��0htOQ��$�ʡMi�뗹��,��d�h)��d�&��v�_Q��66�m���A6�hS�J\��UW�g�"̖q�V�6�9) !�@61l
3��Y-aVc1p���J�*�MV0�¶�вzX l�[X�}��=����x�wܹS���K_�χ��j��|�N�];�q�[���@#�G_Ͽ�'vS��ymP(-��lG��޳��zW��"�cR`��o0�G���*�cC`#��n��N�{սr\�%.����V�8IC�M۲�}1� >r� ��ٶ}�fN�QBa���)^.}��!�YI~�����)A;}����K�$��A윆��M�k�(d1\h�2j���N��L�@�l	����X}o$5&�@C����3
r.W�B.�k싞��(���TW��&G�m�-�����I��!�N�z�BH�%FZ�qćd��Ʋ@�c��f ��D�1ku�zƙ�, �܌lc�/Y���H�l�sJ���Ϯ��,-3i!ju�`��7Zw^�"��{A� �dDT����cE"CARw'#B	���1"(*`�8tB4�# �TN�W�PE	��ga�zK
���_��6;�"��F #o���.3�}q���*Ü���`��.sj�nc0zUL��97-x1WS|�mB7&E�]���>P�>���N�&h���	a�Z�Sx3E'��\B 폈=��֖��Ӵ���i[b*���Uި���X�&j�C����]}Y�p�j(��'�8�h+��U�j�d:R��̂E���Ձ���ٳ�m�w���%S���D� Ff��wn�>���TBFv�F�]�HO�rE8P� ��