BZh91AY&SY/. ߀Px����߰����P�9fpF:��e��	$L&��A6���S��oT�6���U?�
�� 	�&&i�� BD&��mF�4i��@�i� 4�101��&$H�*~�S���y�h�d��z����BC�ҒE�4�$%b@��J7%�?���SelT���q�1!Z0E�=!�Q��rjX��[p�%Lw�g��TN���<3u1�!�]��ִ�HU�t�Y��2?�����uJ�Պ�h����!��g.*��E����G�rHB�px��E�������4�!�6�>�ٳ�~~���/��6�jk�.�m��IA�q��>��s�]��=f��i���aLY�f���S�=Y��s_:�kF^j�m�;6(j �I,����us��)� �E
 �] f���VR)��P��)h�ѭ�;�u�vd���)N-m�]�Ud��d��bB�M3-�� ���V��	0p�N����,�mH���\�~^q�D@�6������a��U�)/N��6�qɃ)�d��d�a�z�f�KSJ��!�+��Di-$�1r0����ȳa�a�W��� ,k���;�����)ێ|ޣֻ$s��O_�Io���>z�/�Β3t��\�xWЦ<sm�|�E3`�5(:��#�D�,�x@x�B�ǭ���q?ɗ6h@����C����.tX�67�����Mi�7ë�tވ%_4��rЯ�9M��<8i�w��r���+�K��.Q̹��5I"�R}�zgv�J�ْ��rr�ee8���KL��q:x��]�����Fs��T�CH		���:��l��P0�dGi�qP�U ��GM��%Ƚx �a�ӷC���(F�����h���-����C�(�02=���xiUM���:���h*�=-ٟaY�@�V���D�1sh�U�a,s��H!e�36m�ߤ��_��)>�6�jb��󅦦I �ҹW8�4;�9^.P��A����^I�X�Ѧ4aD�O�hB�j���(E�e̕'��ˤjJ�.�����QD�{�u"A:+��e3��y F�D�vo�f[계������3w���X`�6�<��Í^�<D#�m<�%\��C�n�F��7��ǀ`�9G�_��-WP��t(�J���1���	�0n�Y�y��d�fS�R��VX:�Eo��l�Hy+nld+`n������'�qp�Y�Y:�k�ie��� 6H�Q��zʱ�L�y�]�k�Y��܌o5�p{�@�Y��b�&'�Sَ.rF��F��sg��H�
���