BZh91AY&SY \�f �߀Px����߰����P�瓽];�l16iJH#MЛS�=�M=G��<���SOQ�z �?D�P    �   $!S����Q�   ��@ h  h�  �#T�3&�2��@d h�2 !� ?x�=`�I/̠cǗڿ�%��QI�`�"�$�0����tĀ��ch�a"�/k��qy�[ 	q�v{1����\�n���Yŕ&7])J2O98.v�H�h*�����������B-Lqc��
ւC6��d'�f�N�Ѓ��		)M��+�xk�G���0lo���Oq��8�c��gڃ�`�۳vo��D"��3�uC邒ڎ�u�h��j�!��"(�w� &�B�X�R�k�rxP�,$���q�֢s��Y�)g-�TZ�q6��WXHa6�"���h�P�_	��3��4�XM-eL)�T*�in�`#p�e��
K��/I3VW$�@��e(�H�*_Y(�0ixI ���¨A	$Q��᜵�� �~C�ب,��W[z���+<�P�y�2���#�B�P�$�5$�����(�	��I$���ľ�y�'��ޱ�Znn�D8۵�����	N$��<h�4��1E3E@I����:g�L/j�$�jر����T��s�M���ƛ[���eן������uN���zp��}X� ���_�;�@���j�G�zs���Y[���xú�Z�`�-+N��!�W����C`%�B�~���8��.^�E*�����tЏAТ�o>��1��ėx	S�KɌl��B=�H����QP��֐���]|�0NT_k\bL��-�f��=�,�!v��v�:�@���F����`@4�	S�|0P�F��%�t�J%�SFd̸�W2�K{�"I�Ŋ[E5��Xg�H����V����h��! ҧ�5�B�����{r�=-���VңCAi�"m���~Pb�N��q�Q�S�{�3�X7(�}]���]�n��-	�$���\���s7Dζ͟�Xz�܊�h<ɢ�h�O8�/�I�RVh@@��]s0qz�p�:�$fF��v3� Ĺq���.	9R���@�u���\�%�J�V:���^�����a�#{�+)QAc5�ss�ݘ�L��!���J�c'��$�[5�`l@I�=T>��Ч&q��3Z�8Ih�� p�,��F �k��#_������L���6�_JF*�-گ
�(o����`%L����J�\Ó�Z4
�W*���M�)
@r[�$Q�h�}%�/�r��@�!�6p,��Z�Rr4g5j���Gi�]V_��ޓgII#KL�������ܑN$ 4��