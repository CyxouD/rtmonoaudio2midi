BZh91AY&SYK� �_�Px����߰����`���� �x��#Z��	�MOSF��4j4bb4441�~@�M���L�����  �     a$ȉ�@ � 4�  �2b`b0#L1&L0D�dLBSz����S�M�(d���h=F�L������.0SDJ �|*-;����G��f��	>�@�~��ࢹ��;`R)xG���z7���
֠�=�`V�����U̷8-������:1����RAۈ�������b��U��nD�\h�q�lAE�?r`�����򑐀�B�PO�3e�@B���貧\/~�4�ʀ){n����0�7�w�2L�����Ն&�%}<���6�`.�81ٖ��2$��u���rE��Bp�]�Q^D�5�LH\�4��˲5i��� x�#��o+a��[+��;`�䲙ʣ��S=�4*^Ғ�t�܇:�kE��34$Ҟ�w'YIh�z�3>i�xj��D?)2��:�d���ž>�g�8XT'�i0����vft$SH�T�p�Fk���ķb������-ۆ���Yq�5520鴊���b6D$�Iīoe�XjMX�	:�ñ�D�`�n56�$D�ف�u�A��5KiFP��ѱgnl�."%�
�I���A5!IVipQVX��ز^�;�D΂�غq#y%C��c�C�OB�Z"�9��S��E�'��_gO�;$�H)`I$�Aa����R �|;	L	�m�!]AI����)6����C��%d��HkZb�1|�,�C�0��HF��48�T�CHig7��	��NUUͣv�gb�K��q��ݼW���>x������3p����z�Y�N*hH_;u��%V�$�K��?50(����<]E��YW�h>�ɖ�Bηq��9�̾��U���IG��%��3S��:>���E*}i���nӖH�nl�Z��9>�$)w%�c��D��������fj� =��+�o M�.�iH�����NE2�%�)B,�=�e��
B�)1"+��JuP�����0�B�-�u�Z�"�5E]��0ݰǰ���B��d�f_=����E����ZE���9kИI	�NN2J�(�,j�yi��}d�mϑI��w����f�pbܖ��ix����0�=�M�nh�}<���]����@�|��*��E���u�:�<ӢV��fN!,���o*8��WyD�Jm0e��V��;*�ٳyQ0��e C#Z�E�k24N�� �L�C9P�.
�8���9�jx��(�O������+���vN�������+.s��r���E8O��9t��9��u����l��BBr����uy�ʍ��J�*��J�B��N���"�3f;5���l�;����a�[[V�Nsd�.}:�E�(�Mp�9����Xz����B���H]����Ә�Nd(�k�K��Z�3���S9[m�J�5K�}ƭN�	!ffGqz����}/f8��,�#+m�*���"�(H%؋��