BZh91AY&SY	I�� �_�Px����߰����`	�}���z   /��妶eQ�$�dѡ�꟢��1O��@�4`	���~CAJ� �    �i����4h  �@ ��I�i�bhhh��&Mi�dR"z�4ѐ � M��#I=!��z�����  h	�+��y[)R �$@(�䘲�x?�
���a�
@DV �2���)/�  3f6�!�Y�nԴ�� Ipzn��ÂM�}Z�U�r��z�фQ`Xaa�a�QAYPPaUe�TXXEXTQF�QVg���wP�M�4�cs6$�ؗQT�Ţ�R�����Z���5�O��(L��c6i$fl�8�P�V��2<\�	�Ԑ��hp���}x�0�$�������w�[�}N�t��la4���@���L"R���Ѕ��m�����Cq~l`ݸ[�*�b�Z/1��Ppw���SEW�Ó�W�M�3���J�Nrǯ���J3M��fa\�#6�c"��5T%d�fߏi3�,
c��T�w�+����!����Hdr#0�$��y��;S��z������_�ƞ�b�]�!�#�R��$x�]!S����h7k��Ʉ*�GN�_MQ��	�du�ﳶ|����"
uBO�I��O���&S!�:�4�Og��3B.���*<�
��/�.�\�gO��H|�Up{n�d�d��s����"��u�{S[\��w
_[�j1����sq_�_#2f���6X�l��(���F���<b�	�W�b�ܮM�ByO\tEVU�]�#c@���B�c��5�N[�10/;�^�q�&(���!�ۍ=��B۝��"Z��(Q ޗ0$��:���I��E��r,�n�m�h��������`'�feN��<4qs��`�m�ډ��;[��GUo/w�9�kgy�m��]tG]H�x��n��F��wE\������@�|;�n*5�2u�NH��旐 �a����D%��V_,���N�.Y��C6"�؎�ddAS�� ^���������[xT�]i�E��߼��������ۢ�������-wGZ�2�N�U�����3�tW\��u�bv̌���Q��H=exc;��e.7]���u���Ar��;��Tr�˻,�K9�:w��]n=�̘�=s=�j�#.̓5xbe�����S������TQ^UUA�	( �rv���)z<|�W)`�6D]���&od�bcldB!��A �a��X�b*��@��`D\@�b���Po��3�5^�k`�&�ٝ�M3czVL'�Fk����9g(6������qxp���l�yN��<Ղ��}�_"xj$������5�w��åd��
=n�������1�@�ڶ~�s��1�	<�h6�"�I�8�3����n[J��[)��';��c%]-�jl?�o�u%�Q�����w��_D��+�'�wRЀ�=�l�ﱜ�]��ы�b�[
v��5��!�_}x��	 �儰F	A�ZR:W3�
r�`u̍�&슍*�"�>ҽ�&/���^�h(0�s��s�6��m�\B
���T�=��kY��(+9�G�*G
�U� 7v�Y��i ]��,2�4�QQ��hq�@}��W��J�u��c�/Y���R'}�͆�kΚ�a��h �	/Gr��F�9L�m�Dcq��[&��meV�`���f�1Bv�UY3쾂DPT�Jp�B;uH�X*+����!�D���s��*�kи`	�m�R5Y^.�(;��^(ixT�G�V��G�����Zb�6�}Z��Z�#`�u<gN��F1I���ڙ.��4�� IB�z�Y��#����T�	l��٬5�b�;M��TzONFT�[���}Xd{h����95�J˖�A�f�Q���%cU�HT9���H��'�qA�V���X�d�p�HxD	�6�@���Ǒ\1^ɳ�i���ޤ�r7bg����sb���H,�hޜA�))zR�a.B���)�JM�