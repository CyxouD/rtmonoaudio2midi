BZh91AY&SY�{x A_�Px����߰����`_z�p�qU�
��D	��I�!�$����������h���MT�4	�*0       sFLL LFi�#ɀF	5$�24�4d    �@sFLL LFi�#ɀF	&���OM)��ڣ�M ��� ��I�0@�H�������� �R
�H)P�&*I��`�1�ta"�*׎����~I@8�p���O���q9�S����75�{�1]����Z*��
#����wmb��6���96�/x��`�5鹸�r�6l����
���,r�: �,m���t����pf�_��L��:�|����VY�6 �ҁ��ǝ��x݃8�tT�U��F��O}��K�/^$rN��6�'����t�/���	ؑ��ikY	�6��\W Q{��5��;�L!�iL�L
����/}O�Ah-���{ʢf;�`�N'$0���x1���Kj�[I�T�����3dSȵz�yA��ӫ�	˾j�Az��YL�5�2���UrD�5*��4��_P�	�x{��$8��BM��v�ٻ����Ajú;ގ���BÙ����&��s�����e��9��J��||j�,��ǧ���9(���UA^��	~b��pv35c7�U�Zq�g'+�֐6��JC��1IE	~HJA`X�e�d�$�!�>W7nP�ajaV��jf�$�`�f���wK�!,���b�A�]���'�2��S���>d��w��Y��)N��PIƮ�>\��O8�DI�����c9��P��>����1�,]86�[�R�*46�Є����x����u�DiM�9��Uy�Ty�I
�˙F-�a��R����ɨ�;��f�I|�czD�5�U��s���I�i�W�eL1�=r�e���_lw�BB��P���]����j͘�{�;'z8��(Y$����ҙ���W�L=��$ޢ�ܨ��<�@\Y��w�Gt�ّ�Vݙ����$�uG
lTٴ&>y��P�Y�T�_qq��sZ�Ňp̙�������nz���$���Llc�'��z����]����ѝ�-�HF�~.k�P��,Ok���b> �E�4�"٩��4ƊH�$ӡ*�B MK�nD�LYFUM:�ԝ}$4&����e�J*�U���y� A
��5��o�&�kI�H��Pv��T(��Eч����������m}�c0v+#�o4��%+�d�l�4�ܞ-:�l� ��G�wq�!��nK��bJ��
����G���7���n��+¬0�\O�j��W��U׺�i"�ryڒ���;q���hd)ZA��Qhхnu37{�EjH-�4�b=���X�g"gT�/}�w崦J�XFzM�`>������-eM}�l��H��$uR;]a?�]��B@Na��