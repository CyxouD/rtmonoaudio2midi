BZh91AY&SY��� ߀Px����߰����P�:lp����� �MA�d<��O)��F�42�4�M4��ԧ� �  4�  %2"I�@�zS@�4 ����a2dɑ��4�# C � @�<�~���OR6Q�F�����	�!�:RH�&� ���H	?�|�G���UM�`�#�5?���ą��ch��EX\קr�ߧ #��w�%�R��U���{/1��Ɉ�Ȉ���'�47-D���ιb�NA!��%��Aj�A�(�I!
��BB1~���q����C2`o+�)�ރ�R��W�mm������Ò𛢕K���J�L߹Sh.�����;�I�ɏD��=F|h�(��j��e�1t��!�%6'^X�g���ǃ�����½��`(IUR:�f�J+@ �+ P#�����p�cP:b"(�R�+��5��R �e��ZL3����:�]�v����N2��x��fʠ���)Y3��tm�6$����I$�@@�M������rz��aV��%M����񬒉@�S-�o�M��`DT1z�Ye'7m�aa��S�[`Ci�0d�|#�u����[2a�޷N{��I~r;�=�E����M�>�csn"�tܢ<3����3ց�F��W¥;x��$:bc%}=���NsW,@��%��D��B�QFC0�@�����c]�e�R��$��a�rЏ"G��+�c���=`"~t�ض��+e	����'\�5�JC�g��fhC�(ȡ���w�5��7;�3�(`�����]1�A*Tb �l| H(Ul��L�\�A���k,ZH9bWfi��[��k�A��[]"I�%$�ЦR/�"�]��Es��h�:`dwPC�%$Q�m
m�m�I�)��π���x�19ޙ��������е[^�i6�"��cc����06�H=�r�f/�Rc���Yk$��wt.��xGK�3��r�L1X:"�4�l��O�i���NįhB�5/}�$"`2��I�3�q�E�M;DQZ$�����3��{
�
�_e�>��#R5���#�id��fb�T��y�<��;�8�c�e4��-�0lQd���k7iJwa�CY�#�2N��4����YT���m������,C�r��ld҂7kĝ7P!�=ێ����`���|�S��Dʃ	e�Ju��3[@Drb��:����9؞��!J�2�<��ղ��.��Y(��+���ŋ�P��&sI�:�h ��I�S��1� �*fGi�K;��c���2E�Cf܁��.�p�!���