BZh91AY&SY�m8 �_�Px����߰����P�:� �qFZ&�I �4F�JzO)���)��FG��5<��T�   �   "" ���    ���&L�20�&�db``$T�OT򞧨i��h�i��  2hEr�o*�AK�)J!�@(Y�{�����������@�b^�y�(H�p*)����u�t��g��g�tϺ��U��bjC��Ƀ�(�i+ܱXg�	]2����&��M�U�K�ԂС��HIQ�$
�q�2���>�f����ӛ�Vv���r�o���m��;�vL���c�跍����MU�.I���AZ���Sf�.(f��:!�Px�*Xv�N��hN�i �#1V���k���F�qqq��V!� (��>`İ|�_虢�ٲ!�dN��Vn,6^�ͪ�:̻Rd�Q�y��Pl�Y�k!�le�T�3MgEHЦ��I�[ќX8Ԫ4u�h���qZ7��$�n�cU�0��nf��B�0�m$ou[�L$H(oN�F[(p�]����u� �[�m��4	AٽyO!)sdߪ���h�,�[l>�u]he�1�Ƅ�,���K�V{� ,^H�9��c����32���9	*�qc_��˼����N{���.��l��8�>���S���yP\o�������u8)�����C�����΁&+���`Q�A���tG��ޱ����GU����կG0sc>a�)���@�R ��È��{C�z�r"�~
����+}�	��tew�VK�1��~ %/$��l�h�u��pilT;��"�rҼjg;�)�;��I�,�)n���g*iV���gU b�CIZ0K5�&K�@4�[�a�
jA`:�#\�=q
�*� $Ϭ�Mɋ�%�\����a�W񋞙�UJ�]��vͮ ټ:���U����("{��Z��F�5*5|��Ѩ�])�j��.�\��� �q"b1ki�@}�4�_�`	F�35�m���#�On��>�1j��
NVI�	v�/xZN����M�ԗ��i1j!���v崑�L,V����h�1�����.)N���]�D툪�$��d �Z�/��Ai��-��03s�9�M@.�
�ޤ��:�a^Q�g�u�lͿhVIE��sk��C0{U,��9�9�$���][��nN ��`f�N^�8J;�	뺳8F��*�|�30�p�,tVF �bkOL!|iț�N��)�RV>1��J�Ӳ���*mj JlQ��Si�E0��-
뫝!~�jmC�1�$���	X6���V,�4B�臭vZ���i�l���AV3#�ң&'�ϭ��z��M��5�.�e�rE8P��m8