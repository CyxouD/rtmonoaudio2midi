BZh91AY&SY�,�� 0_�Px����߰����`	���`9   ��*API�����!�?S(ڞ)�S�f��4��Pj��J� ��h� =4  �L�1�2`� 4a��4�L� с���L��L#dɓ��&	�F�!�D�Bd(���3�$�z�b4h4ѠXT]~���K���
���г�~��/����o@�ނ,jc���uEu�8H��*)�#����e��K��v���p��C�Q�:9��z����K�T�Ȗ�K̬*��*��¬,#,H�0�]�UTTe�@XF�nQqkȆ���!�H4�I�Z,6�l�A�k�}kfa����WE����g*�p��wL�k��1���y�`Q��ʈ�G?q�i�!&``���V8������?��i7��=���=����jf=��e�"��p����S�(�%#y��.�EIʍ���5�"'���q�k�D��j+:!����Li��<`\��v�$&2q�Be^83t�	c����ט��_ �#}O�#�,a�Ie=e3kʲ�$6ezHh��t�O�BhaS�0���4K90�s�R`L�t.�^*lx1)�B�r�l�դ�d.݇7k�I�`ӈ�����[�Hh�A���K^�R�ѼlH�D24��"H�VnВJI�^�{u���aʍ���℔ s���"!�鉒*d�2���ȺǮ7���؋��UfS'e�ڱ��T��Ъ�B�Q���[V��2-d
P�f��ݶ'�zs�t�F�%J�FPh�QȈG�Dȩk�2�z+�U-�beD���K�ql#��+f"�Td�و"%��O�E�"��n�Α�h��f�L��e���Q��%鸆R�؁3I*
2vw�-=�*<����y�V��b�:Z�'����8���[q�-L`����5�Ub�'#����H�r�
Q. =��НJ���Kzh�t��YD[�uy{T���6��hT��q\���>��y�}'۾��P����9*�vW���;bm��i�3�b�T_A:�Q�h��"o%^���#��,����}W:�aT�Wcj�XQx6kצm^�${��6�WW%r�Z�sFN��t;��"6EMN���D�E\���n�pK�WqR�Wz"�#a�u���ݽC�m�\�y���������^߄{�Q_����A$����|KD|�5���3�--VY �������L���UUU��厨.P��jH�Vh"��G�z1��p0@�9y�H|qEdlVōw{��.�r��|3d�v���˚��ן��)�����{v���8\[�^�4K�.���¬��BLU!���Ƃ?��\G��޶U�o_>���DE�_� ����S���D��g.Bk�[���ب|^�o��=GFY7hؽ�0�@}�ځ	K�_�3�4Y:��0j�����o׻axH��~���*����v����[PY<���|"��j9�s�p�B=��B�Q�h��奍���f-i�j=�FFT%�E��g�sڌw�_7�6y�s�6R��+�IE}z!*��x�S� 9�a��E����yh�3�翜.N�b�m/5d�p�Qy,�$N!�[8m��,����4�k��a�����tDs��rF��ݲ��+�|WƂ/�����I�:��ӄ�%�Y:Bd�*!�Xq�����DŊ�]�-�
+Cz1���6e=T�L��:7f*�qV/,Z�E�j��~s0DZr
����ٴ�9PEނ/��0�oSp߄+�����:fn�u�� ���m=y����R��Lγ�ิ"��_J'[J���	΁	9r��(H��'���p���|4����F`f�N�=�"����)�ad.��`��~�R�Ȋ����RY#N4�ǔ鵨@����k�gaR�20��-&J�H]�56�Ә�N�(�m%��d�p~�3�k��T�܌2���%c2<d���i{1��$id��w���]��BB���