BZh91AY&SYk�� �߀Px����߰����P�m����UR	$!����zi�I�����S�&L�� L��`d�di��L�eO$� i�M14  s F	�0M`�L$HM	���4��#S���@�4i�БF܉$J�D@HJ)p�x���|>������`� CP����'�1!^0E�m�CH�Z�k�j� �K�����A7>�:mvء���8�|u��w��dC��i�T�W�MM(8 �tV誦{3\���IS��x���r��N�;�(Ǐ�{�����Z-n
�l��]+�)�&s�$!;���`�0��Jx
T97'D�ulI��\%�m�>�g��#� NJ2�������)���0'3l������fX�Ä�vp����ዣ�`�@��ii�!HTV�@[T҇5g�1M��d5r����v��,�K��aj3U^��4��`���ù���������:��|��I�O9$�@,ykm3�͇��qC�JD9��)�P�����Z��L;S􀢛	�$0��a(�b�aC<'t��©��I�X�� ̄�-SY��Ͱ��QϿ~�\'Z�պ��.�~�=��>O���J�����7��(̢;���x��!�(^��e$�w���%%/\v��Xw��Fů�_�d������"����!����Thl���ԥ|ar�i�c�-�+s�Q���z�D�R�cC@��ң#�$�OZv^�@`�+�9���F	�uM3�:�8�=�5V{'95�yS[=���6)2L.��8I� iΗH�>�C��f�q/?�%�Ґr��<�5\W��m��b6WG��$ޢ���V)�OqOPv��3�Vs��LJKrxET��Yq)q_�$K�tD�H�ՇB�[5�̡�3K�Ω��j�>T�� E4lccR}g�h?+��R�y3v�<d�$.��޼ ���/>g��0�}�芐�c�4[EBY6�4VDbM;	\Ѕj_}q$"`2��I�3��EµMU�bJ�A+I�W��@�T�ʠ�GvH�: G)2�M����4�LL��=,�D<���6VƑ��{�ϳ+f�z7�i����=m�cSh��k�&�]�kn���,��2�P#w6�t�7����ʑ�
qƣ���T����Ep��)Q)�}�Π"�,ę6�jF,�*�i�8��ٝ׾�-��T��,�}9�X.�͓�}(g ��^Rj�T�E�r�6�/��-RL�w`��cC����$f����w$S�	�m��