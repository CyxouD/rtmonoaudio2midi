BZh91AY&SYAp1B y߀Px����߰����P��8tiF��A$�@M�ښ���T{P�(P �?@	J d @�  H�!"?T?T�M�zF�����	���dɓ#	�i�F& �"JjyOS�h���$ 4   �K/����Ċ$!��P$�ϊ�]ߝ�v�:A	�aa~�H砀)#!��u�4��P־����5�V��%��@QӇ���(vj�RA��6��'��	��d�.YA#FÌy��*���*D��I	M5
�qd����&��X=���g���|>�C��8�F�bزk%(z�
��y`�B{B��J�aj�"�9�2U�#��J�G[k�@�Qd��+6�nIv���N��M̲'a)�R�gy�����D��/���!*(R1�`�
(�
�����1�R��ýŪ�@-�h�'5*����ep*�����*Z�2�T��[R["-a�J�Ze�PܮYd$��Zt�c!���E��ޗ�W��g�n���m���km���
&�NҟQ){:�uW�g�fK6DV�kX�`p��#��FƑF}P�m�!�R.M/
��9�ab����͚�I���b�����?qI�_~9��|)��sg�6������?��g���"󍟭X<�垪�������J��LW1���~s%���{"<h�Z���y���t.f6!J��w�p�����*1��B���n�1:�w{�z�z"�}�O�]���;Z��߳%��DΞ ��?4�}�@�����H��=q�]ZD��E���wN�T�we���R�����M�!�p3K����H4�h.4��`�H� ӭq��8���h�*?�H�p��>�Xޘ��|��~�/bv~1s�6b�UԤ����B��0�X��H����L�T9]�8#�m�׿�Ԇ�ė:���‹c�qY����M�1�4����ׄ�6 �ha�a�{d}4�s������͌�W�*52@@���8w.�0r1n6���"�T;�̉�h43�¢e1,��Ɖ�Fe�8� @��u������Jp儻�H�X*+���IG$�A6Q,��y�Br�;�0M����Z����[3���g���}i`t����	�,f��m�p�fC$h�f#fħ�!:�ę'�о�Br�.��g��Se�q�k�4P��Iò�a��֞���f�2(�f�Z~PS�QE��)Z���mEd����T`B���s;�轇'�qp�$���T��Z��:�I���D�^	}����@��l�]���j�F9��`:�!
��u�Ji�G�url�!"��F
�o4)�rE8P�Ap1B