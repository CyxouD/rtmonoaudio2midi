BZh91AY&SYu
� W߀Py����߰����P�97 �q%�%TP$�L�i��d�j��{H��ɔz��A⌏CPjzh �@&� �   �В4�hh4ɦ�     8ɓ&# &L �# C �"�(bh��ѣdjb2h4z�h�.���$)0��@�)��Bx��>� �?ݶ)��w &�����1$�cG;i0�\{뇫6K�|5W��w%N���j�V��6a���2�'b�2'u��u*Y4��ba~[��ƺ'�dV���aK�c��.H$2݃	^dȮ)>d��$�+,�BIVsx�������`	���7|���ם~�����4�m�;X1�����l(!
|Ęۋ�����:)L�q6&�(�,a]�& �
(K�$���x�0�+SN�s�3�A�R6t�΢��/.^�ͻW�$�"��ZK!�4���ZQv�˖-2)�4�`��C�*���P�LB�1-%�u8+,���Q��r�3%�dDY;�YX��E�	��.��վt(��cdp-�dM�'j�1���*�ϫ����:ĐH$�I$�&�rlm�h�!������0;ԈF'zQ����
�h@�����B1 ${Y��0b( �\�*������X�Pa6Q�ڜ���*�qc]���i9UWV��~k�.�,�!=|�]g����:����A��_�N��p�j�����*�BR�3S�
�����Y[�ڿS�I��͝����o_�}��!y�P������nH�����n^��^�d�OD+�uGp��ϖ��b��>�� )u%�Ǟ9��k'I�bz���򴇹j����wg`����d���OIv��i=���n͓��s��u�&I��I��| @&SJ�.M�*KLa+=1�q NYK4ޙ~2��~��e2�qD�y��R�P_>�I�۬[���v������	�}�BXb���)���A{�Ӹ��B��"n��Æ��b�,.��X �>f��G���#�O_�����ծ
M,�K��j�\�a��+M�}�0�| �"�4�Y\K3@�4RD`M;	chI@��]-" 14��99-�H�SPM':*Nz�&J�gy�y���#�����]�� � [��AӖ��C(W�}�����w;�Y�D=�5x��R�H�!G�����Y��'�y!gې\�r�E���%����K:U�<�h�a����4XB �5�~�h�;I�Y�����"��|c;����Bc���v *��.�1}�a���D`�R�A�s,W]�t��cST׎�Ǆ�pn �E�ar^�Ż"4.��5q�V��\��1������2b~\���ps�5�d��;��W�.�p� 8�