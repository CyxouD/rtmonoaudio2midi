BZh91AY&SY_bl �߀Px����߰����`M���y��BT�$��H�ѣM1MOH��Ѵ�hi�� j���&RP   	�  ��G���L	�M�M4b2`����@=M� L�i���挘� ���F	� �(��D��������P�L�@�����)���"�PS
 ���Qi�{_�Q<�+5��H	�(����B^'t
E/(�s=_g7�([�w
E�i��[{�^r%��Ӊ7n�Q
Y�ni��2�9����� ����R6��2�yЩ	�Cy^tu��܆��Uo �h=����?���d�D�.��eٳ��z�����-$ู�2j�5�_.L�Ƙ&��h��RL�D� :m��5���T R�L��h�x�D�n��*�nM�n�`6�f�`iR�E�H����{�Q`��.t�;R�XQgÖ�S2�6;6J"�dU5�Ub�J��i۩�p�W:�j����!֙���f��Ų��'`sA�9��
�q�f45�`����iS̪`�����]��m������) �T�����;͢��̢!�KM��.�&�KX#*e����V��0I�:�iŧ%�p;l\�I'6�<����gg��m'�c��lI6�ޘc&�íE��+*ux��4g/���lp ��P�jo���
b8=]�F]+��x�{
g\�\�q�� m5	�-�B�B���Dk k$ִ��E�gZ�P�}�1 e}'r�����n��h����/��9���Iz8���S�|�!�04'��S����!�����i�$"g\>��d�d$ǛWT��;�-W��Zz{�gf-Iԫ�~!����G�9\I%�f�d���Uy�"Sv'<}nT�p���K�v��ŗ 8��
&>�����o%��LS��[�j���ܦc�E|+g;�!(�;�ye{�S�QG�\��=���1�L{0��JAq"��+S�X��[*�aC�	m�fvjX�h�Q%w��1����7�������'B�f����L�q�/�W?���i��B���=lP�9�X�Yh@n�tE=-y���E�Ƃ�-I�(mA���g�]RRX	�6�����`�|�<�e�C�T�&52-�B:x/P����b���0	�ɉH���x�KԦ�\�Q@h1���D�Xɫ(�Q:,�c������\�P��V��.*%:}8�9z58�0�rN��;zy���6�MLM8q���v����٠:���V��#��r`�	�3�͸�0�p��`��Q(۶�����y���ӆnˠub�]�$Iî�Y	�j��P�H�E�5��킖=��mm[�Xe� ĩs�]�≔Kn�	ɧ-&У\JɁwm�e�q垓�)�EC�H�8�T��N��@�
��+9�Ӵ��3�eFݮ�B(fGqb�V#��kٍ�rE��"��cPe���"�(H/�6 