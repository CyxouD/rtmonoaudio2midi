BZh91AY&SYy��/ �_�Px����߰����P�& �=VX��B	$C &�����2OL��i�iF�d�5O�LD� @ 4   D$Ц��z�h��~�z@ 4 hѡ�101��&$�&�	�x�4�= i�  ��%���$�H���	1H�D���_��t|�T˰l`j~9��\�$c`���a"�1kM�g�^z�KI\|w%�� 6���p<�P�k(4�4�?� �g�ln�T�3eof��YA#�q��3�>�1t �&h��P�w��[�I�7�zb�����/Z.���ʱ�����K����K-9�K�2P\9v40��T�1�ŅQwu���/n�%F.0�g~--e��-P�§�8C^B 'i	m��Y�< �/�#��?��\�mҥ;�[}�B�ݶ*^c�X� W��%�ή`�B1���-�l̋�fl8w�,!V͆9��&x�ų	�`�#R�2i��1!bЙ3M1n��wc�#	l������L-��9L"�n8Ѭ��C�aΐC�e��k���:�`�]H�m��~����I�O���`�%�
�A)z���+է��%�Dc��e��ږ����o�������8y�Z�,L\�,j�����,�]0�)~
��dfH��Z������0��v9O�����2�/��I�����b`*�ל�*�?�	p�?���Qe�b��<����ѓ�Q�}�eoW��\x�35���svN�A�m��˩�q��^c�39zu��5��G2Ɂ�>����f�d�:4k�E��4"~��ޗ&7V4:H��r�뚚�#3�c����v��Q�;UP��:�8��׉z�5-B����g-@�CP�1�0	�l��v�RoT� �;�F��Y��g�M�b��l,]b+�����l�R���= %I�!�r3�:8b�OzpP<2P�8K,v���C�0zXTL���&;�����b��4���tctm2 J5la�a�{^q�s�9��ꖈ�}*��FI��u��t�Vm��>ӘEc�d\��Y(�*'[lcFF�I�N-S��"(X�Jp�B8����T���o4��&I�b��u$�v}4lz+.E�%�	q�� �~�I|��=�k�bz��9�s�'����6�ï1�;���0�1�r�k
pa�J/竐�0�p����@$�.��1�y*�6��-ZU�Vk	0�@p��ȄA�kN�atg��*�:�d�"��|cZ���a@�Fu���T�	J�"4\��QE�9>�Ń@��ڧH]�:�!Ә��%X�\j�iā�/F�r�٘��*w#-�l� J�dwT�b>�{1��$\ɒ/�v�B����)���x