BZh91AY&SY +JX �߀Px����߰����`	~|��P  �XUQ��I ɠ��3)觵5<��6�F��2T���J��A�&4�M&�@h�4d���`F�b0L�`� M*��`6� �a0  �E��CF�    ���Djb���ҞQ�SCM�OPW~�
����r- �� �WŖ#����q�ќ@DQAXa����� �`���x���v5�ֻ<���H]������z�W��r��A��Eq�K�j��D:�"�A-��H����3kP�,��*�&m!V�yn|5��q�Fi~Hc�7<�����h93���(5����	V�@5���?7����I�/�yF뺍��o�@�%��k��c����U�Q�.3���F���H��ɋ��tXsJ	��e塂��4�J.HbwD��,��u:p(�sahi�v���"�k�F(a��q���ɶH��1\6��U�Àh�7�ڊ��R7�ۮFn��6��Ɣ���Y����u�b�9֦E)��J���R���2���p�{���ఛRsAa�q7�o]���1����0 ���犬�`D"@��n�
$�3T�:j+dj�Zw���Q�%���ڂ�XIb���#%l�x�ƌ�M����;"��*`%�7T&��/hF�f$���HY�*�.�L�Y�$�(�V�ma�C�V�d���1
s�����;*�=�tEo�r}��Do������,���E�`��PJǑ���Yx�D*�
�W�kK���Xg��9ɗʚ~v⡉�
ް��A��j��`؜%�����:�@���y⣉�d���r'4�3�º���ͻ��&��q4�VFI)V_F<j-b��~0~k+^��,G�09	�&$��7puI	�9٩V\dkˬkYδ1��eDO;=�ky>�B-��(7P"�'Z�V.����x��0�s
�Fa��j�t]�[��;�l�=b6�<���Of�\TFMx�ͣf�9��ǰ��P=5�4�ޘx�q(y��c3�/+$�[Z�5��-Fǜ��,Ցq[�/`^Q��3`z�:�#4sK����GGI,+dĄ��ʇ}��'x�M�}����Ww3|�ys�x��R;���8tv��1��������<��eHٵZ*��5U�M;�Ts�c͐�Nt����/�����>&����m��0BJ&�=J|�K��|�X�]^��NL�L�A�śI$�Ĥ �8�������� ���-&0�$��,0i���$,�a0ɩ�KX��fH@�b�*k{��|cϟ�͇B�<�xd����)���$����x����9$6��9�m�k��~
rLI1�WD��ӓn��ꘐi�)�a�S�sw�D��^IfY����@�� �ȈPW$"$��Vmǭ�]�����e2x$�=���:Y��v+�1�Q}�%䶱w%�X��aR���"��n�CJao�z�8���K*Qۦ13�i��^'�j�B�+s=�����$A(;[)5��ApvԎ�3ѡa�f� I9�_~�͙��6/�1<y�:D͐�<hS�W��%A5��M�p������ٜ����l9�:���
�J6���%�� �q�Ph�4�����b��ze'E��[a�$	+k�cc�}�������ч;Z�Œ 9��r��Ff�'��s��> �"]�#++�i��6��̀ @��^6"�e��� �d#���%I�"�q4K�d ���sEO@Y5P'��pñY��j
�PU��A�쥂�L��<�|�Hp���vUS�AS5�s]o�P���r8�I>F I5���bFp���HN['��^u�H]]'6~I��KX|�-�f2����~�#�����uW-��
��g�T�k�T�By�Rz�l "Nz���=A[���/����dgQ"��6Y�r��Ek�B���IR'�m��Z��e�=�g�]����9�����ITX�#�Χ�xB����D��2F�hG�.�p� @V��