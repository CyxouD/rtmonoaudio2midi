BZh91AY&SY)��z �_�Px����߰����P;�X�قl�$$�1�52(�F����6��&'�"l�J�       LHEDт=S`�`C9�14L�2da0M4����"H���zT���������0M4`d�Բ i�ޠ�K�J���u�Z����?�W��he@LAX�����"H�8�q��wy�����&KG�ɝtgH�9K51z�9�(f�S��M�-a�����CB[X��,�ʿ�E�Db�H�pĂ1N<$�T_z�F�N"sO�R�ЋT�I$��B��Xn�?#뾔��f�?�z���֊���hab�.ɓl֪�n�R\�H��|F���g#�*�I<�ƺ9'Hˬ@5�' �\�M��,�܆w�,c�ؔ$PZtdP�	�%	1B��H%6�i�T�\{�|'�����	ar�v0��-��M���U=���ꄶZ�8 �;��`S����o6��] Y�LjQj�a�d�udT4�Hlݳ��b�	u�F[ZM��:/���@��VV�L��H�EF��od�����Zn�\*¸T���D]jV������"H$y�$�� 뻭�8�Nm�E��m*��ʕղ@�21 X�T���`�`P	UN��X>(�◙l��&q��m�v(1�M������*e�S*��k����#����砟���>�>���5H���]�?9o�Z�^wm�����I1]c�>��۾Ƅɽl�?#��{�.f5�%�g���)���fbH
�E!%?O0�O�|a��h�J����wi�H�BW��ܿv�=�}~@���/�{o�$d�k�e��	 ��N����yE�o����1�5��?�����o����S"��W ,�a��k�~�1	���v�S8E�+-�c�ɋ�%ȹx�f#_�C���+#]J*���	*�aֲ֍�}Ҏ]	���{Ӄ���ҟJ:c��:����s��D�ArͰ��8�,����@n�@���\i%	�a�a�{d���s���t�����j�fxXjd� ���@��v�V��q���hNA0L��n,�]�m�B1�[������yl,%��m��#�d�@�E�1b��C,6��-%�DBI� ���lxX`����[�Aٿ1p��D���ޔ�;�7{�=��Շ�`�wE;%'�r<+B���NL-(z8��ځ$��G�������gf;�Z�)�
U��W��p�a���φ|3�Ϳ=Oeܳဪ&>�Eo������:l���$�`IF�`4�֠��r|��AuӦ���m#��xH
%��Rv������7_k��R��v99�v����=�Eu�=�i�(g��n�y��7�)����c8Y%���"�(H�w= 