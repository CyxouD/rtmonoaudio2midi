BZh91AY&SY TK� +_�Px����߰����`�M� 	�*ф֥PI �4G�Fh�m&!�4�A�@�?@	D�@  �  i����� �ɑ� 14�0�mI�� ��   ���a2dɑ��4�# C �Bh�e4$�&��)�h�@h�m&�Sv�� :�>`A�,(!@�>5����T��n����@��E�A��@K�D�H��e�'ٻ=X30���P���`�`�T�EY��\)�$:M0��dC�0�~I2yȄK<!�r��Ix���ێ3�*�zE�T���S�(��B�&�
�(�{׽�I�� �Â� f>�Ú��y�ߓR@���Μq�8�V=��'h�	�83��c��mQ��G:LV�el:*)��Hv�h�
�����F�4!��k(�e�	�;�M�o�;v�j��v�;�p�w���(m���u��n��r�//d#��Am=ED�6�%��J3L�J�^,cg�V2�v�JsB�J��V���HTkA)�5+��$S����T��T��U �ٚZNI;e=�@�T�
t ��wJ��
K��jIĶ	Тl��&��^j̹L����Y���T���5#(�bP��!���鬄�d��.��L��`�ՊtDpR灡S�A#�c�`�P��&M��yz�|�Y@�Ƥ`�F[��qk���֙��W��� �Ie��H	$0�Wz��$A<��l2)P+Mv�CbDDԛQ"����R��a�B'\�[B����:R�EH=�.iC�Zc��1`e;�sE�6�l+k�]���S�O5�m���l����s壻|����|�����������|4hRBH�W���M�	$1M#�����o�bMY[֊�΃��"�c$��M��Ռ��Gҙ��"���Q���hvO7з�")Q؜���V�gG�tg�Î��1����Q�EL�5�Cϩ,pF�Nj���j���6��޴��&�8A6н��1�om��S���Y
���u�Eyb���E �
t�P��T��-���alӨ�vh\��j���K�rna�3.�Gԇ_o��Y8L�类gý6˴5hF���w�S�z`a$��88��*FɰSa� 6��s���˗IA�a����4�X�����Y'���`!$F��35�mg�x�#�F�Ti����e��F	RF�E��E�3�o��X3'HL�"����F/R��e��F���TK/2l�l�:�*��S��� b*\!���e�T��S�Ӑ3��S�8�S�9�(m٘�(l�\N�IT�pu�2z
����w�X��S�Q>Ӭ�s�5�EI�Ϥ��e��2b���I�1���K*9/���VrWXb 8v���D f��j3�$e�Lg�gt���vJᆍދe��1*\��YɊ*l��},!�Ң�Xr|��2�ڥ@]}��!���_Br�����u8���3�C�_1}\T����>PH��2�ؕ��q�1��$bɒ4�;����\��.�p�  ���