BZh91AY&SYw� �_�Px����������P��l�GqM���)P�B4�jm&��H�OQ�4Ơb�A����% 2     S$	4�y@�4@4� h��`LM&L�LM2100	B0�<�覧��0Fh�&�*�6��A;	I!9 QHG�ĝ�}�� ����E�$T P�o?L���/"�6���,ak];�7�+� 9����d;��6*�T�4�d��4%��'05G	�S���>i"u�E	SN�'�8�&H��0	�_m��"��$�/�����'��xrE0 �32n?�W��k�
=�/���8��{nT=�[ݛ�*\����ەw��YY�J����J�8�S6d`cVŦZ��8��7	2��P�����(�k�\̗�!�%J(i �%b�Č��IoK��6R&VA���j�����CC�F���jL�T�tY͝�(F3kM�������<W�4���e���7��5$���"I$�@6�l��LG.�b���7dJ8ۭn���vd�(8H*�B:CS����� 1u����pW[U0��v��� �)1[[�푣��U����3�k��v�}︗w��������U���ay���� e����ʬ� jp�Hu�@�|�ڴx��o���+z�.�cg���8ʀ1�[�X�8U����QP����!p�� �ә���WaD�S�Nx���ƹ��	��šy�d�@s�� (ޖ�/�h:tezD�"zmR�I�^#թ7�i�C���r�8�t8�X/��T0J�i�����C!��\H��2iHt��/��C��*�v����ġH ��3L��S%�A��YV��o"���V)��PqL�Ï2#�""�k�L ���AΉ�K�e�><��\CdA�]" ��^Rc�4�b��5�L�Օw�LN M��61�'���}�"Wm�5Q���J<)1�I@��`96��f���^> 芐�c�4[EBY�1��#�E�;� MK�nD�LP�I8wD�2#H�u����6�(֯�� �@�{*	��m3Gx � ��*����b)�	h�=6��A�'&�bOA&k\��va�=�$\B=GA��*Ɍ z_�Й'�ۃ�� �_-���%xcy׿Z^�%�:mYɁ�]����7��NC$��NzX+�8�*#�aRH~�V�+W)��7b��s ,Ĕ���1d)T�̱c��n�]{�m���@r&�=c_h��������3�h�y>B��Ä���hh�=��J�ߞ�$����M#�iY�_�w$S�	 �{�0