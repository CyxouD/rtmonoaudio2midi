BZh91AY&SY|�: �߀Px����߰����P�8�t	�z�K` I��H�<�h��&
z�D�d�4z���J�   � � a)�L�<��� i��4@� h�z��z��4dɡ�ѐh12A��OJ zOS'��4��  �z�*���Ԁ��ER��� s�Zn>/�E��`�� &�4���2�`̀����"���<�����@E���rQ�c%]~Ɇŕ��y�ͳ�*iF�Ό00*\��G5/%
���vI�4�I"�bJ���	�d���N�y��}��y�*���:����h����2`� @����NO�z�j��cQ���<rp��,���j��]��;���D���J�0v�/I4��{r�p��� �F�����&FRf����VO�wl�T01��5U*��≹4��wàe5jb���G1v��w��LB��Ќ[�X�VU6���;�F��R��D�8�0U�փ@QNE光�3�t����d��. n����FSIYR�n![��0n����/iW=�Ws�h>�la#���)��䎲���r���M$$$�I$�D1�n>�O!1�7z�v�dJ77��C��`� w�"��>�+v@U,M�%�B���4g~��a���YK���� L����l>/��~%'e���_�y���La��l Y��2c�n��) �~2�0t���� .����_R����\��ī���ڼ$@��\]��w����+Y���$%�i��| �o�~_L7��%�;0ν�D�m����9�$��On���G��}�9�hƼPE9�%?�^�?�s"�O4e�l�Z�Y�A֚/Ӎ���D�����Lv��1�t��C�[���(!�h�D��
��X��0ʦv��u1	}	�3:sI����kΘ�Y>��Fa���~��f�XUej����d��yE�>�}'�R`d�Z���Χ��[���Im�5]:���A�+Gy#�ͤ9���y��W��	J�&�6�����|��cZ���Vid;B/���Ңu�3�8�h�ɬ&	�H�$^���IPZG�P�N*" d(�[� " 1"�	��tc$��E6y(NN<�T�hi��!'R˶`�WE��!-BǤ��t�9Fݲ�wޖ�}�OĠ��vه�C0o\L��:<���m�*E��l��И�8����I�]S��/����r�k:V���
�bI8���F@�lǟ)�8J��`�].="�Ld*�Hc^jQ��٢���*�j�%F���k$ͮ�$^èLs0�*W�m+뱶J	�ᴊEW��
廘���c:�/�'z��ѯ������3#�kR��x� �owH�d�\?��]��BA���