BZh91AY&SY,��T �߀Px����߰����P�8� f(��5�BI��#4��e�"�Sb��4=`LM&L�LM21001"��0�C	M7�!��B49�14L�2da0M4����"H�I��i6��4ѐ���ʮn�H��*��Q��G��?߆�	?b,j��C�p�@L!"r���2ǋK�ѵ�@���q\2?�g��5�8�.[��9���FC	�2���rK�L�$�̧��th�}P�f$0E� ��Q����7�2�{Y���Le�W�6�ј7���\X"�]K1��{:������i���ps�c��s�{h���S��M�qLp@�"�q��0	���u�)��+|l�gm_[-��q{�RFq���OV����m�Y�'d�B��X�*���g�a�l�)�'&��[���+'����R�P6*���K���y���ɶJ3#�C��ݵj��0�u�/k�f)�VR�Z�S'Ytp��vR��'A:Y��\om��;�5Jkm�,�N/c!!U��~�<㔒	�I$�@1!�}�|�G��%E��O*W!���7{:�61زU8����HZH�!�Հ��&G=;�:)�X��X�afH��X���w���NVY�g�M�������	��o�����x�^�U:�����([��Jb�߯�̷&T��qk���^u���b<h�Z�����i��7T]�o{G8s�=��)���A�R �忀�㩵�,�D�r��!���q�h�S�F��ϩ���!)x����U�D�'Iޑ����(�wd�"�g�~�3�ǈ����t���O9~�m߳{�4�;�M�T
��E؀��  �1�B{�XZ��4?��F����g�b���(�� ����=3d,*����E�2x�^�޷��qc����B�(��A�=iP��b���XDn�H�֞�7ُ.�Ð�n$M��p����Ih�41%s0�0�=�Ϸ 7lG>��d�X�֪<+9YB�ֹ�٤�C�1�5�R\3�&DŨ��a���m�L,V����X�1�N:	p��pPs(ʈ��7J���
@A٫Cnb�
-8���2�78s�SlE�-}JH7��PP�v�>���9�ݙ]%9͎v��ҫd�A���S�!&���D�'gw8`�BNQ�S�;�Ic}��cb�+C�j��a����Z��F �q5�Y�c^�li���
S�VZ>1��J��
�cʍ���Jl!(�t3��g�Ea��^4
�)l�3�ch9�	$䶐H��`���m� f��c8�}5����с�S��		^̏#B����mV��6STb���&���rE8P�,��T