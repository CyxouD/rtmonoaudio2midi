BZh91AY&SY.~� y߀Px����߰����P�9fp;N)�٠���A=�6Q2bmQ�zS�2z�4<�馠�=��	(L!��d`M��@h`JdH��4�OPjP  @ 2d�b`ɂd ф``(�(i�4=&F��4�4M[Yͼ��,Q����AgI�`����sd/� 'P#@�腔�t� H	t$M�)������˜�n�̔/�aJ�@��:���a��@�B
!	$�=�f��d�kI�M(�Dm�4��T��%
�ˉ���1���)��l�UQa� ��q˫���`Bf<|i�oY�ʻ�����1���ɸ���p�29�X�:UN�6��RH�,���.ˤZ�zձ�@%	
���<}ʵ�7)��iw��,N�W�s��^�U�k�Z��K�`�q�Q
.d�GfK�D*�"����+"��Y��LL�`b��ȶB�DaŔK A8J�I��aj���v@��E��XFd��2X@��]���vy%����\-�3�.f˔����uF��GĠF�D��/(����}��$$$���H�B�m�k�Uy}[-o�ӹ��(�ݲ��&j���Rr40.��<PhD��i �
���F�����B��s@���m�f�
Hi��>�z�:�N�4_�;�MGo�6�Oo��Ϗ��������^z~�7:�t�.�0B�������_�LR�˫�/	���"<h�X��;�r�o�s1�ZV��veM�����@G�Q	(�����O[BX�r�>4�]�9�1Ѫ�My/A�8�i�_1L�m�h2t���	�'����bC=�_��s�\D^����9�A���������6P�Yu��b��3�PD�Օ �Zד��̂[�8L�F%�[cPFW1v�2�^t/b�7��Lي��*�W���G�c�[�񼥆8&Bޜ��:�є�R�`@n�D7�=-VӫOCI-dN!��Pq��Vj���`!F�,36w�'��|G>��,i>�;�2��CHp!u�.�39���Kd�r �%�yH���~l.n-�#�T�r�`W,@
k�AQ,�5e�Nݪd!fݣ70�@�����������vGv��k��@!k,yʐte��P�q�>�������iV��w9�p���fu[$j���$�X@Fk˱�²���7kh�ߺ�<ʵ�Cf�cE�-:��梖�f�N��q��> ��wZ[�l���T�,��R�5�&<����@�6(�l0�(��'�8�hW�d��WF�:s$�ȂD�^{^���!L3��Frn�J�R���cn��G��m�}5k��(���7�He���"�(H?C 