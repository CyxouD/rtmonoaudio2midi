BZh91AY&SY[�r /߀px����߰����`^}�l      a�a���i	$h���M14�H���{Th�C�L4� *Q���&M0�C����0&&�	�&L�&	���`LM&L�LM2100���54�=A�����4��D�$�4�)��OS&��Mi�=&�=Aj�U*��YR��P$�i ,�����*d��C���I�#P<���p@��'l
�I����[�0�a!$jzij����F��(�jW�/�����_�ែ>���Zj*2"I!�i�dr"��V"R�B<�Kr���f�ӤɆY�e)�)e1aԔ�9�%�%���Oښ�d�<��!�s7�e�:l��-��L%�&��F��g'�.�� Ԉ��F	!��T��"�3X������ި0$�Р�\�.`1�����B���|u	^�u��&�I�k��:��q���*9_�`A���>\�{��V�T�7|���/�h?���M6qrl�˭�ٽ�gL��T���V�&��B �d�@�d;�.�b���l��?
�Xm2�4��߹.q���mD3714FS`h0�;��<��KF�SsX�a#i�j����,b�BM<���v�f�������>�����~Uw�=�x�e$��X�:�T
���}6'��[C��.GB��u�<�R,��Db&·ğf��b���C������*CH7�_^t���CaA_)�5k٧W���4����H{�vF� ��6�@dk%�R(����a_ �bA��H��Sza�ǩO�	Т"!��r��7,���p�aP���LYcJx�EZ'H�!�(*LHa(u\�$�{�	EHYFB.����(�8u!�a�D�0/W�P�Tn�U&�"6X�(Xp�ǌ#!DdG4��.dW��3��!`�=�M�k�:�)�W0�1^�w��T�I��F��m=�f��B��A"u�h���1��]M�;Z��d_4I�J-@�{7p�=�ݎ=@�4g*X��-�s��YZ,���xR�JDq=P�7PЁQ��
<�8Q���rB������{V8�*3mk���	�N�;aD�oH����Z�y�������kܒ���S�+�����J!��A*#�L�qr}X�RN�t&����^���+�ؠ�;�ZU͈�d����VW��vF���\����rhe�ԭCv�z�̙�A�C��b�5I9ӳ�۽��9<��(�/pq�ŵU���1Hf�@�H��JևTU�]�5��%��\���S>���N�7��`�ǝQ�j2��dL�;Uꋸ19G�x-"�u�$�����[ߎw�����Ȣ+�J"�#7hB[}uv*m&�F��j����yW=tj](�Z;��G��a,Z�A�|�짢��楬ң�A�[�b�7p��]U�5u��s�����+d@� |"�|��!��|�(j��2~�2�P4�Jk�:�kճ�w�GU�o`���C
���Ti��w�ցd>ً�Ν���Ә����Ж�At���۳�-�����u��+�f�o<��wƋ�v�24���|M`c ;��N��V�\gZ�55�����/�`���τ��k`��6-u_5q5B�1"���k���O���>�$I<rI$��Eϛ�����~�NN/���W�!xz3[CH�xAT�qd@*J�����)DF����6�`QRdh��N�0��9z�8s��	"�-b�����O�Iֽ������<�������[�|��M~�f^[�W�f]�͊�BH�߷�����Hb����dG�w���ik�U|N���P� �QR㣇b� �f1�&�RP����!''8�q�׸��:Ӆ���d�4&B����'��s�@��{E1�?����K��Y���Ϝl�׷v�ȋjyu{�%W׼].�V�b��ۧ!�ώ9��Z��$������� E��y#h�R��Z-�3,���z/�0h�5�FJ,�$$�}������~r���0�����l
��ک���!!$T�=�b+��t�>���k4,&�'�\�y�q�C��i��.��%�F������#��7l���Ռo5�BH��fl^�G�H7(�}��lӲ8�� zE=^w�����S�mg�
��(��A��$�C�4�[˳�E ۻ�	p=�fjݔ�ᒛV�%d��EX(�mZ�a�($��m�d�v�t�(�X�H�Ě���з|C�������p��	�-f��l��m��hd�#����aR0��+z�����ì1�HIQ��s��ꜵn�V	iɳmV1;n�d"t͉븺�{h�nT��6�V���r��h*Hۮ�́EM`��{�]�ڻ�|)�
7���KVU�����po �-�k����4�:���A�х��TV9�6lp{ �F�D��X�����i��N��8m+��6��H�
�t.@