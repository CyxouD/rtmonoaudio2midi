BZh91AY&SY��@W _�Px����߰����`?z���s����$��CI����<���A�L����=L�Pjyi% C@ =@2  hɉ�	���0 �`�0�)�!O"� h  i��2b`b0#L1&L0H�@M
��1LSe�4d2z�@1��ϰbEPE���$�G{~0��6�P� b� :C�x>I �`�1�z�CH����]��x�@�6�!|�
Ԗ�+ʩ3�D3�s:]� L�f!�PYӲ�3�t�;�M?�
�$��"�� Fmn�=�ں܁\O�c��]�ԃPU���iI!d/n��=�L�``�x��}�M~�{Q��ȴ�dە����w��K���1��ü��!ǘi�`�Q4_i����5"�l�Ё�� '�mnw~��p/aCQ�ۨC�tդ�9iL(J�H5TP���E�Vx-�s�8gL	+1��%ܧ�t4+g������GT�C!�jT
�E�p��Dc0�`��H�sZ
 ��wl�I�� j��Eִ�#2�w�f`��Vq�����mK�Lj�:@�;���zV�0\��6a��9m�'�VC��/#��W
�d�$V'l����^I		-�I�"�f�d3d��6�S�.�"��s
S5"��
�J���i�d�4��P�Fq@FY�Ґ]�L.^�~m�o`�I,���5�g|��SO�&,9N����c�~늻��f������TK	}j���*� 7a����S�� 1M#�cv~��gW���4��Ο�K��Ȯ���6��9|��f@������57�?�]b'J��珹�A��<,�͝�9r�6��wܗ����CSQdq�������r�+鍜�D�2w<���(�W�ȴ��;'!�k��y���ZƐ(��ZR:V�1����w�eJ��@��o�3L������>���޳�ନ��]�K�`�̏��ܷ&@*���R�s��m�aA��)��)nȼ���i��o�T���G��v���� �|Llc�/��u�R'_�q��9d�����ڀ_��@����<�'0�#��.!��H�ʪ�5�1��#QD�'$����Б�/R�<�j���TW8������l�Y�ܽe� B�G/U���͈ڀ ��.A��i��ʕg�=>5�1D���O[������nlA�0��̑��{O��+�� _=��<%����X>� B���Ƿ�.�&�T�h�!��U��PG�JT"��g��n���Ľ�\/��(���E��5�j˝/�.$��=N� ���fSz{�UF��7j-4��f�1|��B�9�$`�ܶ��✳�&1�j쥜�5w�+PQr2Xvv@y�@���ޫs/����g|BG[M#�c����ܑN$<x��