BZh91AY&SY�$C� �߀Px����������`�mp b�R
�	$�4�Q���=Lɩ��ꆘ����JP Ѡi��4 SĊ������h@�!�  ���a2dɑ��4�# C�	���dɓ#	�i�F& �HT�3F�~�解MM�)�=F�G�����G?��*8AK�(Er_]���'�P|~X6�0$�PcP>�� w܈��H�*)��͵����ʨ�ʪ��#�cэ��K42�C��!�"zf"a6�M5Y��JPQ���738M�p�$�J �a�`�\~����2g�s(�U��&r����H�_z�VaІ�a4K���#��<7{��L��00e��,�Gջ�CQ��~�x2˃p��p�gF��Sϸ�:*�	-�(/�$�B\oA�N���T�ZQP�P��@�&�\�-QN9sM�I;ҋZ��7�������@��<��)���z,$'��\+����Lr�yRi ui��|���i�.� $&�P�e���Yk	LJp���[�4�8%�&�A%L\�&n�4�+ .y$�M%�!s1��?Q���oz��m!&���ǜփZ&2���ؗligi`Sl?�-��T^L+d�x�z�eu,0A��6��h����,j��@Lp8��9�yO�WAV4�a�Ka�˃1:�`*z���!�O���{����3\�/`����;y+u6GS��7tvL��_�w���k�Ol�I �[�;n����}���}�uXB�窾�L�`PxD�u%�
�0�hQ���祻�@T8�V*��F�:n�-: b��7�����2HW\����w����N�]9��x�<�_��g-�������r�ٕ.�ۋι��%D�.U�����.� !qqu�+l	�#�wӾ'(���[n�̎�}
� �Î���1� �)�L��$�������z�םm�Obъ$�}i����q�>��*�׵}�5t ;��x��S�\XוF��'MH��=va[�@a�Zh����w��R	�W�o}��i0�Ƅ��k��$Þ�P  ZZ9D�9mx2hF�.��oq hڎ��+Ȍ"/Is�%����O�U܃�%o�C���-%m�J�ܨ:�z]�d���L/�k`@��Z�)�GL�Թ���C����\P�~a���6`��(�c=9�SP���fl�n��&�ʶ��[��t6��_:��s>�7�5�\�\�-IpfN@��%D85&W���F1�\���Ļ8�1��-��\/46e;�6ަ�ɹ�U�ť�X(�Z�/Q�4�ǻf�V�Rp��At��Aٳ9QCl.���0�1e�����d��pUM�״�9�qN"�����k���V�n�GRa��p��kIr�K��3��S^��Fՙ+�}!���i���z�:�q�7X�~T���N��+��R�Mp�EE���`ڦ�c$�K��X������0�ku,ڬ������pp �+�ט½o�9��wZ�A���STr4�l���@+�dr4��~�-!�Sdb��%n����H�
��z@