BZh91AY&SYz�[� �_�Px����߰����`�� wR��I$���BcI����d���2h=��EP�@�`F�h hɉ�	���0 �`�0���H�ި����   �挘� ���F	� �"@F�)�T�G�I����Q�J$�ݶ�%3	���!/i��������~�Te�6�&����)/j$��"�m!�Y�v�.�=YhB����@�=b�K��^+`7dI��h��a�2(6�r"&���tۡ9�Q6�MOmEX5F�BBd��}d�"�wIMB��x�*ըB-M]Qj���,<Pf
��B-mR�d/� 뷇��قh���O�Ό������5�]����w��+�:]�u�)���R�*s�|0a�S*���<��`\Yh莏7Vfj�-l:�<Bmb-r0�E��qO��Ft9�W�6�d��"5;���p��W�.�\��U��.I��n�5���F]������:~!����S�D[����-R�L�/gZ�
�C�q@�4�{"�X��\�d�_q��ųDc�F;�l��.dBV^��iŤ�N�¦RӴ�.vi�����Y�!�Q�V�S��n2��9<Jd���.#f��9�������i\<;	�NK6@z���m}�f215f8�6��`���!�6��5�L��FQr-X��'�lU	cA�1�1,ƌ�cSW;*�X�r��/:�� �%%&�6�ܧ��ۻ���,�\E�,�3{�7@.�
bĪ�?XK�H�y��Bb�¦x8:;腓�5/�,��	�
X��������OEqWy�sNu�a�{{������oǇg������!�r7�Р���>�^E�!	����V		��%�w���w�/ZxGy�p��jl��-���G�yݵ�ȕ����\ frǸM[~��Y0�T�oN��#�9�dy�|��g�z�f�@u� B��-�[�T��#t�Wh�>���H�-l�zq��?�K
(ߞ���3��۫�q5j��Ml��+	h%��H�:��iҸI� �L��du��UjP!9�[�Rf�K�������^��)�FE��YP_�ҁ��N�G�$E�ѱ0b�T�Cj��"�'(P}�
p�%-����i���3�.�Rъ��.��H�3�Z��*��cc�|����H�|�+��̴�brL �f�^]ˀae����@�}@ꋐ�qk(�*�N��4^H�Q;��p;�W�d��������Fa`���*��EHA6Q,�w^���(U��&�\Lhȁ
�Wm'AͣX����J�>��:`_��j/Ak��e�F`֠�#q�k�+�'͗X#zd����X?�)��$�_|�Pte�-
ĩ�XBVxv;���PsVo���%���
�S��E���L�֚��.dX��C�tX�V�4�F�V�L4�U.A�t,��͆!�n9>R0���E&�٬�Ej�y��Άr5ZMR�A�˄���AY���mU�0��sKf���f�G>r>�����)�֢ߨ