BZh91AY&SY �h _�px����߰����`	�}��x   ��U�lZ��$�&M	��L�꟔1M�2$Q�24O
�@F�2hɦ LCSƪ��F����41�2da �i��s F	�0M`�L"R����S��M��C�2�b 4�&�DA!�<��zG��@Ѧ�� �@�B �F"$ '  *AgQ��"��g��S���iSP��K)TH@F�G+i`�.Y�O�koBI.�����c����w�ɩ%7r�ҋphFk��\N��x����JX� %n6�e"�-Q5"+$t�6�lUIhӶXB9)�i�+�:69AX+��V
�$V\��C)U���j��6��?K(����wќ����+�^C�V��=�3��� u�)A���C�ܻ��<BJ�I�VM��aݭ��M��W/6���@����6����0�C��p���aG��{�1Ǐ%L���UW��n�ᬢ2�~;��B?���9�o���_e�9�:����V�6��7
���e�J?�bA�Ɩ�kd��� �뀠�+!|��T� q� �j6��i�D�HY$}:�/���?Q��Y�	�Q����,уJ.��,�NԑǏ��� Q�D��׺�7u�a���o��AM��TW��T��<4��45u!�N�:��O���K���-qMo!�/H�M9#����,i�Be8���<C#�}4�C�8�8�B���CB�kp��#0�@�N�o%��ӗr9@ZvQs�$w^�&��m�'�z*�i,u�y��T�Eds�:���8�xT�܌��*0�L0�D�q	���<�a¤,����9��
7S�p�ɞ�;��^��l��6�|�j�l���Q��v����_#�vf�ʺ�%��fl�S<z)\ɹ�a�긐��������;n�m���ʜ�a�aR]�[�.U��'�2��_�؆)�A��?DA�^.,��0�'DSd&!��tS13T>֢���G��	�V�ŭ�����c�{l�coY9A��A�z&2ni���n�n�m�CXo)��Q���O�6�n�XF�^S���qb\Zz��ݳ7=�C^�^j��ɥ ��X? ȉ� �B��/���؊�X{v��i�.��ؽ��J���}�����=�F3��uâ+Hth���=����R���ۈ�/9�83Q��WdH��n���ۥg�c�P�6��k�~����}�H$���l�IA�ɱOA)zvxj�Jς"̖rDV�i*���Ā�Ć�����@)�B6�\��I�&1BI&.f1����,.�`�y֗���	*�X���w�;=���̳���/e��/���(y��������ƿ�1y�1w_*�TBI/,�_��W6�$�a��q� K�Dz�_=4jU�}�a�?NZ�d.W+��� �}���ʕ�x�"�|� fr��&����������z�sGYLuxt]{�Cz����U�俈]a;ű��mzDu���_jQ�kᥜ���)�;��X��c����}��j�v��K7R��C5�KB�` �#�	�k�L���`�m�fGp�t�*VJI9Ķ�	�2�4-^Ta��nع�1i+h�����$�����x�GV�)���I�[�H�#��R�`@of������{ui�Z?HТc?q#p��:z >���g�cX��Q�f������ϧ��m�c�\���05X]@/EWӼ����t��	��"��|`ꋐ�o�FU'xi��9��N�2�����H� ʙ� �\#�������Ĩ"��D�}�s�U��)���fn+�ʊ�Ȫ���6�������}gP����	�*͋��1�����)�(��F�X�U�dЉ��)AӠ3lBI'(��x}5�i��.��+��1�P#�V%*@o9��pSEp���n17Q^{�&T*:r����E�7����$��!$���Q`�r}��Ɓ%���kk�����Q"؏^�?������WFW8s�%z�M��1�k��I\3#�d�c�s�{1��R��3YL7'�]��B@�Š