BZh91AY&SY�ħ J߀Px����߰����`O�-�9� �UT��M��i��b���S#M�4�@�ɓjy	��        9�#� �&���0F&bH� ɠ�hC@  �0L@0	�h�h`ba""h�4�=�����ڞPi����H)�rIXH�HrBD�8I���_����YQ��l`5=�)/��j"�6�,!�\���z��f�`@�*���df�S�kv��[��)}�d��t2�ĵ(2`
 �H�ї2ʗ%�f�|Z0^`U���U[�A_EE�(0�|d�1�f_��\�H@V�H��B������$���图��y�_`j��]n�f� ]�@k`��F�!�T����J�|�V��'��Ȅ�*cC~2 '�Ť����!���;�EkAF)���$1kՊ��o6�I�����Lk!�Ҩ}��e���ŹI�D;��HY�Le<�l��8���aVu���,$0wԜiFY��ʇ�Z���K�,�3}8��4���B��3�)TVd��Ȋ� HA�y�!�':/����9jm��Pe���ѡn�ҳ,�SH^FI�5`��BX`��Q���Gu�V��3�A*�ᨺ3Lb�>�߇�0A ���I  AV��x���ǆ�\��Q�)R�~� � $��! C<�?���b�1|�*e�"��2ad����}M$�`�f,ɰv;�S�%=4���f��m��݂�Q�|
�]�����v�����S�����S�H[3����U~d���� G�$�8�z&4�=qS�l6��ks� A�[��$>{���؋SC` ����_/��F��mk��)�(�-r�rN�!Ѝ�<9ט�<�,�h��c����/�t��zD�	�u�� K[�^�g��%}v�kLಿq��e�lҭBުh�u `����7���-)�k|��j��`wb��QϬ�X  s�v퉛0-�f�� �c-�Ħ���`�T_X0+غy��u��Ș4&W	�er}�xx0���r<�,��b��-����}�Aa�*|�5�P��9-��ҹ��W�lc�_A�r�ԉ�Ǯ�����,�09ZHG8<{�����Q��9�P5���zE�U'A�4ZH̢w�Bj}�̑�/R�=Ў��`+��UZ$��d ��K6�/ap�*�p�`OwfF�� �p8���5��X(f�\s�7��|���jz
��9ͿOaڶ��B�v])ZX�@���B;gL��l� r�>�BGG�,�T]��<jV��w੠62�A<��E�g���M����]*θ/IQ�"��~zliI�KL3P+"h��d�0]�Ї�[�!M�5���<� �%�å!�8$#X�`�V�� [��r��#yN��c�]s��V3#y�M;����������єq�5��H�
 �x��