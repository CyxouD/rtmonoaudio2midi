BZh91AY&SY��. _�Px����߰����P��l�N⌴YbFHFA=M	⚞�Ѧ�F��OT�6�����?@&�P4d�ѐb	��0��H�MF�z��S�6��4�L��	���dɓ#	�i�F& �"@�x������P�z��B  � �F^MH�)	I]P$�������LŃ`��jr�&���"�m�!�Y��mش������\��%�� )֭.��P�k\`�xb�30D8�3L&F�H�W�D�v��IC4Vl�q��_|�01%�a��m^t�]�HHV��"�w�i���צI�!�<��W�<OM˯s�ύ���~�ml�nu뗯md�v��(� ���^��ɳ��7p^�87�M�C����� �FHB��4;�������҂���!��Cp�2�qmN��Xw[JX�ĹJD�j�&�W�kdC�J�1��
SТg6̦h�0j��Z<$[�	� �+���d5��Z�6caa��m�#K�])��#3�4�E;y��C�I�O#m���"'7mN�R����cV�(�,�|1��KD��JsP9p}!YK
���"D�!��:ݲ��.j�ne{$��5�w�ߤ�Ȕk��~��?U�<��脹�`Y��z?�V?��$λ?��y	�tխHB=��}�~Es�!8���Ӯ�>���e�w�<j--z�W��?��6p�#RӞ]A�g��p���G���5�[z��3D����!��R�7�c�����aj�.B|�����C0�d�[�(�O]����=��/㙜�)A;u���R�W���/�u楨CÊ���P0,%�W��#��N�y2���*6�\ņ�ґg�S|���i5��D�b6wP�l�e5ԩP_��yN���uȍ��q�&!���Z�䌩�S~�~�T�������1 ]�sl+9�B�Ʈ�`�f�5l����ᢌ� �Qfv��G�P7u�W�W.�6tZ����7Zb��B8๖�;0��2��W(D���!���LW��:c1�8JOr4��MO=RDP�u)�3�߲FA]R�Ŗ1*��UQ&jv^"�B!P#gM�>.�&�i�b��Et6�Κ���+�GG'iOAc5�scv��0nZY#P�q:�M�(0��ٵ�L=�.��p6"�F�_I��#�����QZΕ���7���J�N$�0o#��k��]�s5݉뚵��M^`Eծ*˒�M���3�'Q�E��f��4M�'�q�h���T_Um��HxE'D)�l.K�Z��@��*��6p��3RU9\k���A!�dx�*"ļ�����������_���)��p�