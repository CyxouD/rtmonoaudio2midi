BZh91AY&SY�#� �_�Px����߰����P�瓼�p !��2LI�SL�m&���Q�jO@
*  � �   i���#LL�C&h@ѦLj�4  4      $�1)��j=M��4��:5� 1v�!'��M g�������e6]�`���P¢��q��V6���(��v�-�[1��d�֔"?�8b�璡�2�FR�E�B'���t������N���GxI!m%6�HgD�͎?� �Ǒ����J��A�*�$������b/,����q���0m07�l�Y�P]����I�ˁkje�D�r����//��+��מ�3J-+���L"m9� tN�:�b#r� �A���%�vqk��1�!'�H�ː��,��$��+5��%�
fD�!c
�.���AQ �r��q1���ua��J�B.S�����x�rc�6$-���8N@"�@G-o0�)�J�]Y�A��]�	�[E)T���ywE�||�mF`��	�.��ms>�.Z�ݲf`�6HZ�	I�����=�}_�(�A ��I$� ���U��L�}�dibE��VI�����ǃ������C�n%��ť��`$��¦pxNj��&j�B��`�#,������/lq���)޺c[wx?%n�����?;�N_.���!|��G"�	n�7���S����t@�t����&4׋�Yi�m>�R+f,@�%�Uu�\[�/r$��%�93������R�}J_;�C��ˢ�1�F�\���c"�[ J;R�ŕ�N��"l�z�����=��%���v�bR�v����U���[-����������Ў�rh�hAvI� iΘ��pO�
��(�0=��)$NY�3^�&������_�"I��%q�UM> %�O��D~�#����@���;I;��x*����D�W	%�"����1%�s[~��P�Oxs�L�ke�iMg���61�'��:��D���S���K\�����e��GC��w>NP��#����	���T�����ɧbX�  MK�m��LP��p�aj$`+��8��IA%Uf�e��%
��,	��fh��%�Yn"���%�C4/g�=~��EA�A��ؓ�Tͅ�k0���0\��9#�<�v�J/a�I�m:�)���͠8��')�'|��29*����]rZ%�s�O@ld��9n̝&�>��	��]�]7��L-~TD�Z欹Ϫ�S�,5>,	WQ9���kF�B��5eV�y_ ӆ�$^��@s&�\��C&/�B��&b���r��OZ�������� J��S�,K~�is�,d�jwN ��.�p�!�G�