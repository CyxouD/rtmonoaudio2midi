BZh91AY&SYǣu ߀Px����߰����`�{wy����T
(��OhQ驴i4b�4�4i���h�h�2�b�d�� ��M$��4�d dCA� ��*i�OP�&� =FA���挘� ���F	� �$LDJ~�h	��6SCG�4��=Lf�����I ,ĉ��
��������U6Y�`� �jz���LHA��ch�a"�.k�z��ӆ  :���I��s�sS��V��[`��*S�h$6�2�%�&������	)It$;�<K�$^l��ijQ4'
�TO�d�m��)�E�n[wtC�i�R��dF�Y�O��Wt�+V�1����<�Θ��z||�b�쇓��p���p/]�|4Ê7A��J�߈�X�1:����p��)B�U�:�̘�mp��	g���uOir���M;l/p8��W@\M�Y_%��޳EY��h��m;aڑ(�GB�dX�e�U
�ƹR�4+Ei�\a����\�S��։TH%%&2����ȭ��[5}^C.0�ef��tT�q8�i5�؜H����/F��\I�1&�IK"�bZ����-�Έ��nte[S�g�\n�1�S�:/!���9;��K[�k�m��(;����F>�:�c˴ĭ�$d��Q��r򢒍K)E�l{�
�V�8��\rǞ^�.&llq{�;ԩY��3��[s��f�l�`a{$�����]��3-W�a��	(W�Wy�uu3jvu�f��ja�QxN�ck��N�5���:�@k�Any��-<�@����Y����T
IGo�8�����*�=�_����/ d�N]�n�ֳ�dXzvDBp�)1�x����k]�W`�j��q^oo>�Z� �� D%	&��l߉�I/��u�Iu�U�gdE*T����؂lm1�5��X���rI� �2c8�/1����(X��asT�V��!��N�V��D�v�M;����{�4�g#6}�ʿ>8x�Fn���LXW��؜��B���8-�e4��D���]���R��Eh�Y���eց¸=6��}��b֋á���������[VK*T|�"G$U���R�zvt/�f�PE�xz%��f#��QT]�r�+���	�`�λq8C��Jy9+�hƅ��F]v��>NM@7�u8�8 Zܜ��i�#�	Nt�F��=�T0F��� D�@9h+˥3;�w�4ep��&����U5������� ��Do�֮�4��@JJă�N�m��(L}�D��	%Š��9���%	�~�8�� j�B7ճe�-�`�X��;b���h��-3�f�U�Y�o���Bp<��{��kfY�s�"a�{��!���&���K�i��I�RW�!	�|m�!�.RN��#u/�j�(�iMA%Ug��* @B�GG��>n�MH��wid���>�ծP���z��9��%7l �V���H�AgI�ϛ�c ��G��GRe�xp�;k*�m�����L��]�-!V2�Ax9	�"`�g��'��m����b|f�v�	��]Z⬷^���2�=�>K �����Dɷ�z���A��Ug���\���H��A` 7H�#���[��8g�|0p�o�>b٩�FkK��wH�|m��Y�?Y�٣db�sM"J�s���ܑN$1���@