BZh91AY&SY�)-� �߀Px����߰����P��;���bi I ��'�h��l���)�S�f���G�=4���� 44� �@ �BMS�=2�4 4hh�� � �`�2��H�bJ!�(ze=M �4 P���}$��"�@��I�'�r������S0��F��0����!^0D��<, �$�ָ�-��߈�۳BY���po�uWQÉQFMl�b��"J�SR��oXٛ�D�5D��}:X�k��p<b���*���#�D=�zBcsĄV.��n����$�!�07��:uj�{n_�����mY)��N����C�z����ѰZua�'�ɪ�q�( D��2>��7PX�L>�ҥ4����Z�v�n�����"	[�yJ�Z�0���p��]��:kB�u�c;��vRX@9m�^�,䇝TԦ!p$�S������\�'�)8Z��%�Fh�E����j��Gp�;F�J� ܠ�L���V�M��3[llm�m� �o��S�%/_���i�vK8�-{�Z��#���)6�%�B_ɢ���b�!��a%�K S(,PakR���i �3+k�n��~�S�O���w���}m����/?g������������+�S�Hxٳ�����zP�2Qo����~�4j*zƟԉ�e�_K�h@���++Z?p�.aP646?0l�9��8ߟ���E*9)����7���=�6�Q���yz@E:R�����r*�(�qH�lQ^Ec�C�XI|�����%('{�w���X7�&�a�p3M�Z�ިP᥁�]v
d�-)���L뀈�%�q��\�����I�fw�*�*1���(E7�y;�SV/�0��(l�,_�ۧϷ������ZThD�gSg��;$��Ն]e&RW��5�dn`���VυѰ� �Օ�a������ϣ���/�cZ��
NfIP�u�k���E'ŦA��`��n�,R�u6�4^H�);��B	����"(X�Jp�t쑠Y*OX�PE"	��f���!� �{'�{�.E�# ��N��]傆0�dC���%Pq���������9�]ۈ���#0�y��GX���=XmB7&E�]����=@!�~�>Gw�>�)/�үJ��%�6�0�Rp�y�!v���ÿ_1$�^�d>PS����:�;�V��~��if���-`"X�f�4�Idh@�vU���]{�B�H��p�H���\���m� e��ʖr�,�Ob����q�S���̏:��K�.����,�#�â��rE8P��)-�