BZh91AY&SY�(� �߀Px����߰����P��[u�*��!+��"z )��Sh��<���S��d���4�%	���` d��0���=C�h��z@�  2z�挘� ���F	� �"L�G�M6��iM�z�bP=IBF_T�,Ċ$�!!,�"Q�|��?�D��8������� ���Gsia�]}K�fZ �yU�ģ��Uq][Z��3����ܳ�����mUJO�%Ϳ����B���QD��}Z��,����$c�e��׷r�g��!^�$HD��8gų���0ff77���߸�β��rɊ���6u���3T��rmE�f��My��;�!j��V��" șU�Y�ԧ������$In�%�TL�}-b�i�,��N(i�u��P]^f�4n��$!�,
���1P�� � ��hF��3@7��AW��ZJʓ����"vh��@��g%�*�lXt�Z�C7���3/�ua+�p��fh��m��7���A�I		/RI$�@@�M�\Q>rb=:��0�N��G#v���%L�Cd�4A�"*�͊�s.�Y��H/�-L.0���Co<$b5j�6��ݲC�I	��u�t�\:��|/ጟ�����]����$��}'��i�2�p�;��|I����#��7F<���IK�|���B�b�ȱ���<H^�`��l�~�<η��?ű���9��U��GG
��s�A�\����"�$����:5G4�W�R�j�rHr���h��JI����Ya�+o2�9V�H-���:��5؈��l��
��M)����H�1:�*4�Ԁ�:�n֙�����A��[.�(���"�b���;@F%v��QsO�B"��Ƙ4�P0�r)��ܭ��2�$OK$䀵[�JZ]���������W�������0�X�����1ϗ�LsI��'U818�H^P�� k�q>��ǽ�"����!��H�EBv1��F��84!@����H� ʘ)N�G5R1
��*��B\�!�D��w^��B�F��wi�����Foi�-*XE>x�צ�V%�:�4ow"z
\��hm�f���2F�I�:W�0&˗��L����~@��/���i��<R�Ҙ4AT��I8v�E: �����R1 _J0+'�T���)��Z�p�Xߞ��#+�:n!��Q�������z��6��'�FJ��E�&ԼVk?9���fr)��J��Ⱥ���� E��\��q�+َw9#+&H�@�v��w$S�		�M�