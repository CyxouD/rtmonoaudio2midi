BZh91AY&SY�ƈ  ?߀Px����߰����`?��㔨 ��	$# ���H�M�<)�@xI���244mA�~@MQ@   �   ?Ѫ�  4     �~���ꘀ4h   � �	���dɓ#	�i�F& �"!5=S�FI��1L����M4�J|���Y�IP��z@�ܾ` �|��}ʬ��`� ��a�@�4��ch�a"�/k�5��Ɏ�p�^��
:s���e7J�R�:�.a�$��P�	!�����	 o��<@	�dd�	SN�8�,0�Fb��N�Zf������B��!,E�q���>=7�``���qд�]�nƓ_`-�87aso��c��[��Z0LSUY�El�w�����2r*��k�r�U�;C<�vf8�*��J�>�̨�w�z
�o���w;8�wE����/ts'D��%�K� >�-;R%�-"7���Oϩ�ec3�M�C��E�+ Nt��X��.�nX��kb���/E͂�)�3,	sr�#�t��E�g:AY&�kk:Ѷړ5Z���L;e��r��Y/�r��ɕG��2|�[�c���g$dڦF��h���hP�6[A�R#%�y��&ah�	��I ��.
���x"R���*�)`�;".d���f�/�-��7@(;Z
5���(�@i��^*i���ݪ.L/j�����@3"�*b�������Q��_���k�'Ww&8K��]�_���	�U}(��,*�FU v�����Se�3I5aB���q�xԑ�A�WF>�a����1�{/Ű6I�}����E������Z���55��K��N�����\Q�:h�ϻ���Ѐ����I��:��#|�Wp����JD����g;n�)A;Mq��B�\�-Q9#Mt���ޚ���H"��s1)�<�H4�\$�H)���:����J�H�-��3,����b�2��bS|�%��YP_߀0+��tGT��m�6&	�q!�R�p��m�m�Q�$���)r�/��׼ĝc��x�7���z�r]�:�n A]��ǜ����¤N���{8hY@`l�Ig8=}������|�(��Qq�2�����4Ƌ���'bphB ]�l��8fH� ˌT� �(G�h��WD�"��D�c�z�B�GO�����&�r�����(:r�,3B�����U�F���OA���6}\ñk�BF�Q'�vqɊ�1����:�0�p�gA����|��7WI�ݷ��,���,��62�A5�)P�yw�B٥��*�U�(e� �|�����'),p�S�p0` ���6ಔ�&J���B�,�_�g�^�/������=ف�*�mXZ��g ��fR6)*�=�\�@��=��[��|�u�$oi�p�ن?���)�F4@ 