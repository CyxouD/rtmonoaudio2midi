BZh91AY&SY�9C @߀Px����߰����`_-�.8T
�Wf�$�d	6�~��S�M1�d14��4i�jm�U4&� �@4i� hɉ�	���0 �`�0���D��@  �� ��2b`b0#L1&L0H�!M<�ORze4= ��=G��P�e�ܒAf$Q$	BBF	>�%G�` �~���v�*���̤@��$#!�,����E�`�5���e�7�{�K?� 0t�m�#��nb�o
U��$c����rȄۑ�2&s ��L6L4/����b9��J�+����v�je��IMFP�����HY˔����	d.3�yw�Z ���/9�d�mұ��N���dq ���n�򛷴4Y@��}|4[�rY��k���
���$��-�]�ڶ�uHC�Ȝ]�E��%��Q,F�Q�	E&2��BK��KJ�X���)S����΂N4��С�D�WC{h�ҒR�N!TLِLaaܚ�(4�r��Y1�
�ȩ�4�x�i��i�"e9�I�ӇY�h�Sli�aM�e�6Bعl���̭�Ĭ�H�L�U�ڈr��YQH2��$n0�VFC�"�.A*���Y��SU���f^٢��5���ry�xP �4 �m͹O�%/��몹K�舻%�.L��͋c"M�%G�H�����'I1��M0zi�L �Nr�4�L�T1C��WvA�H>y��[VS�ny��'�;y�?�b�?�^T@����"6<��k� A�_�?�.E�!PETђ��I�E�$"4:ZJ{�Z)�7�&U�s�� �b�����	����J��B�y�������\�H�X�J$�hUt���t��^M+�cd��@��1}#Ff�Y�]��ݣNI%�\���=�"XQGn��g�S>�w�$�Z�?�����} `� �ik �;%� ӭq�E �^�.��dp̨ҫR:Km֙ŉ~�R�A��[/x���l�VT^^  Į����F��B:0��t��A2��`�UqE�έϴ(?O1N�$�P@�o&.�4jޢB��4e���[�MF�����=r�O�(>��8��k���Ш��&12HE� �ط�S��ƙͭ��r#	�����Qz*�i��3(�����5>��H� ʘ)N��GER1
��*��EHA6Q,�w^������Mv�Kh.]c�l�iP���N�HP04qv
��gVa�=�$sGQ�~�,(��GX#�2\���h!K��<�������:�*\
�V�͆��"n^��n���@3�:��k�P�]�ҙ+�L���Xߎ��� ŀ��꣪��*�S!M�3-Z�a�q��'��0$.QD�i%�z�W�I�;�vr��}J
g#���=�@�6��6*ݘ|97Kg���4��$z����w$S�	 ��0