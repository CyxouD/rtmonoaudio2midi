BZh91AY&SY��Ǯ 	�_�Px����߰����`�#pr� ��" ��$�dML�M&�F�
3SF�yCjmA�~�R��#M�M42 hd2�2b`b0#L1&L0j~�RJ M @�hɉ�	���0 �`�0�I�@�zj4򞧔��&���� )�4ׅ�A��8�9AL
GA}����U��Wm`H	�j��aT>"#�1���E1��{y_���������Z�L:<���LZ���PK��ӣ	�T@������
�u#ۅ�Y\Q���H���p�6`�M��mX(P ���c�le����\߾��:iE�k��q�Zwc�������6�Ȋ�n�׏q�ٛ� l���;��CB���%`����ٌ[S��g��{�믷���a��JSM�^�LF��O4쪜��������Dcn{����' ]��DU���UD1^��L,0������4�ۍ�۬Mu2٪��d�(T��Y �=�i����@��`��ԡ5��s,�)�#P�L�,��^����e�7W�YP���wKA*�#ȸ0���8�i��yg&�dI�X�U���7��H�����m��hj&2.�H�4�>i%�uL�Pȓ���Lso�r�A*磶v^tJ�vG����6/f��W
<���C�"���W�NVP��z��4E�j��;n�ajc��F�q���h���T�FWJ�Eq��%� ��A�Ӄ�/3P�ʆ��.�.�� `�6K2��ދ��o�ؚ�ى������NFU.[7������n��T�f�!s,�P���v�V���ύV��Nh �ȃb-������p���f9:��Q���x�w-�Ƭ�^�mw0�"bH�[q/s���������^�Z�������r5'����M*�2Tsqջn�lK���#�G�T��Sγ�vLGmZv���I�/�۸����{�]a�����`���IA�)��Xj���O�J̛N��sW'ҡ5f]���H���9�pp�f	ʨ��{_j�������]` :� $$ N>��I�P��{���B����0�8H{�C�E|��c��
��R��(�l��?J�&�&�VJ���@��G�
2�N�2 g��Ht@U$d6Cl��vy{Iʪ�tr[��]�����a眯���|��=>��R-+�Օ�D�7S�Z�$������+��K��>�`Q���V߿|G��W�|M���2�c ,��r`)7��#�uD�P�	)�����O��pK�����oY�${����ӵ��@w�I ��/Vf=��%��.���	`'����'�h����JpN�d��Ҭ�)��YIC4 �NCQ���aDP��9�U�:����a�F!/�v�K�o*-�ǟ{�z�r�Cx�U�8��٫�wǊ�:���1�Z������� �=��y�F�sQ�Q�P@n��v�=+�&�6%&cL'q����@}�,�]KĐ
5�a�a�{m?L�ݱ*�{;o�~�t�c���
#���<@�I��OL閤�5'PK�ED8��sa+����#C}�n,& B�m�A�N������*�`�صhr̟����t�~�������*�<ꀵ�$��B�CW�!���N�������+.s�M�q�z���#�s�vZd�	����L=�.mۃ��	ʎ�>���K�6B��,�Z��J���E'�=�"t͔�FX�`�L�>pR�1%c�l't�C�l��%�*}�y�TW>��|)�E����~��h���t�<$��i�,���V��йx��A�]��Z��r/�թ��Fdy��ɉ�f���;���&H���w_���)���=p