BZh91AY&SY���� �_�Px���������P�9m�'sN�)'	$��i3S��M��52i�F�d�"�L�C&F��C �i�L��C1 "�L چ�h��  h`LM&L�LM2100	&BOBF��dɣ  4�$c��I"�H�H� ]�%g�@Go��,���!�a��).�	�*����EX^׋}l�ю@#�Uvj��4�)�oXJ�*� rP� e�Д[D�Y_��9�A/p=�"��R
�*1�	���f̢��̃ ���B�YP�i&��<uI0f�t���m�,�*<^\�H��0a���U�P*P#���6yX�ĭ�<"� ǥ��mI��Э�earp����fhȋ�a{��z7at�*P��F�#�e߅�,�vELf���mEƤ[,�X5�jэ�)�60FUk@]2l�¾Ps��q�B8Ƈi!��gRƗ�.q�9BYw��������Қ\T΂�
���S��_��Ϸ�8	 �I��I$ @A_�~`�=�T�M"U!��J���\�rIHD񰁅͘�,�FmLX4�X\����,0����K�i � 0� �+r�2�K�N�>Z@w�����z�Z;|j����U�7NW��*@#�f������j1L��Qn��k��烦���U}��������BfYz�Z$:,���B��������/�MY��Q�Ȳ�D�G�9��Y��C�>=��^�:P$� D��mcEc@���#K�#�'��V�T�o�={�-�DE���x�o�:��{�40�u䦖uR�8iXh�
dᖔ�N믓5;Ď�rXs#����\1H��+�Bf�q��B�2��7"SzJオ������pO�E��q0h2��	aE��M5�k��1�OK5D�nɠ��]����cfz`>��{���#W�k��(6��}�#L���J<(32HZ G6���FV����(�`;�b$��T'H�+$dQ:�{B	���"DP\^�8uB7�H�W�+8�M���&B	��f۲�* C�A�{'�l�� E�#O:�r
B�Q�7T�y�]�����9��݀����HGI�:5�icwG�2\���hxr��m���%~:��B��*C�u`E� ��a�@�:�.�8�L_*��)�EAP�
�%e��o`$��,�"�.�ʚ�q�r3�؃!Ъϟ5�ެ1{�_y!d�6H����/�k� pB��K9�Yɱ)Ԝ����>0@�ّ�\�;�����9"�L���ܖ�krE8P�����