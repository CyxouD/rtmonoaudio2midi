BZh91AY&SYf�\- M_�Px����߰����P��ۀ��N�:c4�I$�ySڙ<�=Fj��ɂ4�����RH �@    "	4j�H�P��F�1�=@9�#� �&���0F&$�4Q�M0��bz��   	B?䐬Ċ$�H��I��� �~vTe�6� ��?�@uPI+��G[iac[���9.� �Ilٜ�>�@M�G1NWeTEd���@9�ci�cm��v����M��#/l����`����F��*2��:���R���I"�qNqk�<7��3���hѰ���f�>���z���l��^=;wP�1����dEn	Pv��P~�qx����q0��"�iN-��ëY�v�o#�c��3�N�J.���,͈b����ŵXQ%h]�i�ijC�b�YHi�.�֬�S����7:�3I����se8iO�U�r�Cɶ�$���3	0�3������� �f5b�/{���#�k:9q���1������g.�_��6���#m���M�{�}����j��+:�,�f���kY�"0fg3��kh `Q��b�J7���&�
�p��3�0j�kK�Fw��6N�sJ;IF�>W[f*�������������>~�ެE��<����U��Ԁ]�|���,� �qC���y��{��8
JfXQ��vD���3�Ulj�"�A�!p�������nw��#{�j�\��ڱL���+5�G��G�}+�cr���@z���}c@����&H��L�v�JCə]%ϙ����,�9΀�\ѽ���J�%���h�CF(d1+��bS&�iH4�\$ƐS�A��t�\E
@� ',%s^�}���������H�o!q[�US_� 
ҝAϤZ����gי0h)(�%�N�l�u\�Bc��O���]I _��Pe�o��0o��j�8ݒ��L=�61��9���}.�����,��$�0��.�2B9Y���B&`:��4I�N��-$dQ;�BJ���"DPT�Jp�uꑘX*'x��Ĩ"��l�Y���
��+�wj�ȋ@�
�yZX'��t�=>��1=A�s{k��ނ��9��X��Rd�Ñ�j8���d���e��#��'ݴ2�� �S�؎O9꠶�!Bƕ!�J�ca�$���P���9�9s>�O�&
�ʳ��2�����J*�[�а�SU��@�S)�!�k�{!K1̪��6Zs[s�E�	@k&�\C�ȗ��i�e~@�C9��#b�����n�:�U�#��P��ˢfcS����$aS�����ܑN$�W@