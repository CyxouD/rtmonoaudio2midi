BZh91AY&SYL+�� _�Px���������`�&�@�U��I!1�5<�2i�<�*`�44�4�S�4
J�#���Ѧ�4����a2dɑ��4�# C ��T`�&�0 �0L�0 `LM&L�LM2100	#I��4FQ�<����G�ѧ��h/������ IM��!C��*BI8I��%�����U�0laMC��DҀ d0E��;CH��ַxoe��.iU�,�`�����ǅ�q�U ���4˂(��d%�ޑ,( �L �x�� �,��&N�5�ˋ��j����lq��X��y�fg���;�{iwr�$Z�H �������=9�L@�00xj�U�>�ǣ�mo�v4�U��[�ׯ)P��m�9Tw�ezf���/@�d�b��6b2��VQt�o0�a_cq&��v0)�*`��	r	�H��1���H �#v��q�Z��CuP�8G�2�ie�ة�8>�@VE䚠WB:*�N�qmU�b��
f��N����ܐ��L���ؕ�)�����{6@��&"3n� *O�J��M(�v��2�p&|{����\�� Be�$]cɐ��Ȟ���-!Q��������{�2@<��.(��N�v,�cq��'
M��{%��يK�:��4��O Қf�m�:׃GC�R�XCC�sa<&�Ow92u�ᲖZ�5�����;�rr���0����l��y�DO9�b�$!lV�$�K����M'�M)��f-n.��������þ[{m� J&�>�>(���κ���Z�LE�,�3{ �IU�c���� @�SDUpy��6�aL^�4����-.�`�{�l�����ر��w�r�'*�᧒ݧ�n���˺/���������H���M�<�tS�L@�}�߮�U��b�������n���@񨬭���_q�p��*.f2H�/'��Ͽ�8��?��2���	z���]�h����ܴZ�%?j��CC��o�<B9�pڿcu�8�� J}�lc,�@����W�]E�5��ܴR�*g;��JpN�R{�VOA�D�iC;��NC�_��>��	h���A�$t�2h����:N�%F�Z�Nk#�ɋi%��g��ц%_��=3\TF�TT、,J��7"#�$r[n��|��4�+Y@d�1P�#����C���i��/.�:������37���'J޾�u�q��c���?� }�"q��Xv�sЙ�C�� �%�Ի ��g�#��s�d>puE���DaURu�1��F��؜ZI%j�$E eL� ���T�E�����Ĩ"��D�c��,$	B��w{���4�Ѿ KZ�Q$X�-5¾j���N�������`�Cz���a��[G�:m�,(� I��j�0�p����r��/����6T]�o%�-ii��������3+@�z�.S_D�͂�ga�)�T���cb���*"k�7���b��ЇqZ����������:B�4���Ǆ�r6H��ax*ųi</]u3�k�o)+T�.F���|���0TI�����c�sޑ�&H�c��EܑN$
��