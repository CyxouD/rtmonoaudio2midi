BZh91AY&SY0r�� a߀Px����߰����`_-�q�T(T	$)�	��3T��F���P��&�d�5= %H �     sFLL LFi�#ɀFO�DMM�@�    �@sFLL LFi�#ɀF	��"���?SQ�=�oT� �G�����#.�,Ċ $�I#!�%g�)=}�R�0l萁�a���$b0E��80��f5�r��:��!�J���i���"���A�kkeC�L� �N؝�]UNd����튁\�[������}�Y"/�t��!Q^�!������fS3YZ�� �,�r$������n�5Q��<���!00g����f�@����t�Ձ�!�s�|��vn�[�k\3�lG�4��iڍ�}aR�)4�n�ǐ��A�	Ӿ�E)uW�8's9nշw[	enR�$>jt�6��MSSmD=.袲mi)F`ڪ�]l��*I�[y����,۬)D��F3��94�K�Q�R)̌�\u�J��z$-�%rB��K>:�L
�iR�[:;��%�=J�0p�C�+L7i�^48�&Ҩ!D�	xut�.�Ck!T����Q�V	&�*$M��93�}�fS������ii�k���&Q�.�,\F��t�]��y�� :@ HJRI����IO։K��調K-J�1vK;�0���A� +�@ù���b��a%-6��b�\Ui���|�9\a�U�kk{2EL�b������Q��~6k>�lw�`|su�*���|�{{���%�]��y�%z�r�B�3�xx�h$qK�ߜ
;(/l���v@u��g���6��Y��.�b����8����B�
ὡ��p��y�9[�O2Ɂ���9��{ʹ#�t(��.���r��zB�Iw��Ӑ�f�]�"�E+���$@{,�]8��ݸJPN�1{櫖B��h�)-B��kg� `��4�!|��>YiH4�\$Ɛ{+�%�ۑ�N܊�
�R9�[n��Z���e�����b[
ʋ��!���_H���;on����eu�gPYU颊8Br�!�$��TH6��N._���3'�;7P�+U��뙴HA^Nf61��|y���������\��9�!#�!�x�#���;�S�E��.CA���ª��m�h���D�N�D	��/�"(*`�8yB7U#@�TWqU7�("B	��g3��X�B:�\���kG*B�=�Ƞٗ	`��h��YT)w�z
��s�-��`�X�#�o8��,aJ2B�V�Ga��qOPZ�!�"�����I�<&�%�v�i�,�U(#w.�C�5Q���Ǭ��Ұꂌ�^ʇ������C��L�k$ �� �S���R3d)�C�e�|�L0�-p�HxE'�	V5֥�\\dP�h���N�.#b����iu��A|fGa¯E�w���c[����$g�v�B����)���50