BZh91AY&SY�,�( _߀Px����߰����`/�5� �4B!P!$Bb�MS�{S)��joS�#5=@hh5OѠ%T��i�  dbi�� ���`�Q�2h��10� ���&L�20�&�db``9�14L�2da0M4����$D
hQ�OF�T�Jzh��� 1=I��$����I)����!T��9��	/���0��E�I5?���@f6�Kia��n[�u��L�vm%�� (��O#�89�J���?�Pj`0����$�t��U�Re!����$睧=a�3U��c����($fu�'��%�^=���c���{] E��Z����ˢ��I3���6͜O'���7���҃��@OI���V8p�v8��J�͛�OTa�Œ�rMr1r0UV,�m4���װB���H�]���tљL�C۠���%��c�i�=p����N��ˣ�*��&qJs�،��14�pŠf�*�Ҭ�Zu�F)I�խ��N�;�x�t	�]F\ͳ|��v��g��S�7W��ƣnf&���3'��Z��!dM]Ī��V��k7X�1~
b1�"�Y�_
ˎe�A�U�R�S�@;��[�1��ir�cٙ�'�Ur�[�����%n���Ѫ�DQ�!�c:��^���'�q�"/)6�;�{��'�Njr��ײ�n�쮖�uW�Cs�xw(��ǀ�U�0U/r7E<-}��S��$X���qY�f�D�O~�I��e8"�*���x7q�v�]������3��DV>U��3A������~�����|�	��%���IA��ҧ�%/���UzVyDY����!a]�%�d�,�)�@68bP5�Ш׵�M���"�$��0h�����4�FR��:�@�2E��sc���'�qΪ����,"���������0 �a����zk�P����a���K����@±,�^��)V��m��^-3�{�΁%�^m��3o �!x#���_7���v�u��&�U)v�!:_�p�<G����r�iր��_x	*w��1�k�i�<Ѳ	�4��J=�܈��u�W�3;��%H��]9����'��:Ψ��ΐ0�iC����N @4�\I��S�\��dy���	(���L՘��Զw��1����%7�ȶY��?P	,�x��du�'�������%J(0�:��F�d���$7^D�*K+��e��f!�4V�q#h��:wD��<��X�	)[��a����svHxW��Y���ֵa ��d��\zװW�#��s�d=�ꋨh5���P�cLh����v'��W�H� ʘR�;auH�,*'x��ĔrL�e͎��X@��u`�����t#`	-�$��*h8m�`(퍻�oޖ��_B�jH.1wn~����4�)��Oį,`$�V\��NE�]=�P	'^�8N39x����_�-�Z�%pp�� �1w[��%}�l~�dq�wт피�EN��*����r��U�P��}om3%V%e��C��̤�u	�^4K[J�:k��� ��"�e�e�J��"h�!ݙ���^���Ӝթ��	+���iR���uKg�)M4������H�
�� 