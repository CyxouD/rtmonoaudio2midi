BZh91AY&SY�MRW N_�Px���������`?��@�:�CA% I��e(�i=M5=Lh�z��OI�F!����S���U!�0   	����a2dɑ��4�# C �$Sڔ�A��A����44  9�14L�2da0M4����$DM�h�'�<�2M�I�6���@h��4��?gВA�(��!#�9���_ |��R�6�P���R _
	��1�zXCH��-}=K�ղ��@m;aæ��P������23-X��saK��㩍��qj����<���½���fv�&Y,�zPjE^����\		\^Vv��E0�_���u���̓s�h��(,����å!OC�\���Tj�ňe�|y�.�9�6Ĥ��:h���h1r�V��MzzPN�K�VF����f�1-s�&���Ρ��\��6�t�5of��"��ٽXW��A"!�9Bp�a"���T��"C��x,��ݘ�|�\ �EK�N�f�>X`(�����k���%@32��X�`�,d��`o��ezx�^�B�B���h��̗3��3�iZ��W�p�,������Sm�60mg6���i��i�������*�1jƆ/�����������m��4 �p��S�J^�î���ؕ����6�!�,Š�����c��$Q���*ٜŀ@����i��1j�Y��m	&ĵ3S)j�o��Hχ�k��6��<�I>O�G��|��]��ߺ���ڶ���}�t�@A�i����/��{��*xLK���r��5%2/��:���q�� �Y�3� k�y�֡N�� �:g^��jM��ԬĉR��<��n�t�s��yg��2��c������Խ��t5�#�R+�R������n��,x�4I�+t��Mn/�g��^e���Sk=���C4��H[��斔�N��K�-xI`xjGYsϬ�X  s��퉛2-��z�k�/����\��,Ǹ��p�����Ç2`� �\$7�.u\�4֩�� 7E�:�J��鯐�V[^�S�c��WM	�l��mt7  ��F61헼�r���eo�s7�TZHds4���w�hB9_]�/{�E��TX��i"�����4ƋI�'brhB MO�m	@S)�3��FB�QY�T�h��'�#��& u(?.��5��*E` ����t_Y�(r���߲4����H���v���(�둤r����pJ���0#�2\�0l�Xq����Kn�s�}2[�y�
��IǾ��J f���YR��,c�'t�Qdj'�-x��X�~Z< A�s�G�F몣FB�k�j� �n�q$,��R	R5�P�ޝsf qB��:�	��.�q28|��,��-R��|��Fc;�E̙"�G�0��ܑN$-�T��