BZh91AY&SYv��� 5߀px����߰����P�9lp��L�Z`�I �bLi=&��(���g��������=	=I &�     � �$6�z���j ɐ �9�#� �&���0F&DF���C&�M12z�HѠ �@����n�6�J�! �"�I�h�W��{X-	֊C0��+25Qt	|	�aK�0�����v4l"�TvZIG��2U׭WR��5e�*�Rxf���?9(S�J(H������8�H���2)�i���nd2K�] Ⲣ�G�Ί�y�d$33����N�=篱|��7[I�ځ��Q���[6�LS��Re������	��ƥe�a�X�'�h(��l�8/�X<�T5P�e�y��(�FzY{��L3�*�hX`a&5���4[e*!��P���&� �@��V*B-�)`esX�h�RT�P!���!
@�&e�0YhXyWi%R�)��ty�8���D�歅lLK�r��;��I�1w�)R^Nֵ�i�����mI		.d�I" c&�q>�b9y��/J���F��X-v5Й�$���K�AX>P�!�*M�H]p9I��lK��	2��`�3!"��V�sw�)����v{�p;Wd����-?�
���W�ч���c!¯ڋ�{m+�N*HH�_ן�S��$1E,<��s�����<h�T������=�9���_��C������)�C2=& �|>Q��8��vsJ���]�v����X�n�5��ƋYx!"~优�X�,d����'���)r�%��g;�!)A;}s����1���a}�5P�+n�M�b#��#E@#�AB�q�*2�`��&G�IQDU'�!�Y6�S�O��e� ���=3ZRM���V�S�N����B>�����)FC�zС$l�:�>�f!�$�0�TP�6^��)P���1�1���`>�t��M#U�35�mG۠�#�G�4˵�Z�LZ��ۍ�X[�?u��jSr3��IJ��8�.Kj$��(N����{�!X�C!D��IA*4bBl��b85b�76�2MBJ^� ً<��-�<>;����"��H���f�̂��U�!����A�F�Nʫ�
˜���C0u)2G@�{��iN�	�;P�釳��hZ���3�=���+��6�ҭJ�ꒅ��1�;�!v15��]5`�	X|৖���C�V�Y(S6�CɌh��E0�R�9�coCrg��&�/s�N��襴����85�H���\���k�@��rVi&�N��g�ӥ��+fG3:��K���ns�0d���g���.�p� ��_�