BZh91AY&SY�Kk4 2_�Px����߰����P�8���SmBl�8I ���i=M��M4����j���de �    �B!�h�  i�9�&& &#4���d�#J!���~��cDC��4Q�Lng���.B��쨴�|_�)�����@��R4���]J.Qq &�9�R)���n���c����hD??i ���޶����*-�W�+TJ!Q�H!N5MP�#�qS��Aө$&ȘF�i}M��9��i�Ʊh4���>B�"��+�TSh}Y�V�&��E$$���zY�w��з4+�^I�Z���۳�3k����L>#8r�/�/���84���GW:-�e�PɎ-:B��5���I
�M�&��)pl�z�f9ƖXy̷��u�5Mԝh��0��\b�B֨��3���"C��O"�����+tH3d/kQe���d�#(6��Q�[���F�F{,�֢�Z�	Y0�d��q5��QlE�3�ʨ��j�A3j��~ήn���	�"I$�@�b_ɺg0��n���8��{��sD�PA@63Q!�@@���@� H���A"$�9.�m4v�Y��7�p݊��Q�1kc�w�r�'+,��E�O�#��`�n��S���|�|����L���L^z�]�^�4$ya�����SHa�A����Dz�e��y��Z[�Ar��t�����$�kWkXk���aGΙ��$���Q����o�bՂ"�~)����Y�$z�����wl���'℉y������N��0g�����$(��Gն����E�5�fu�68��X�rȰI��p�]B-!H�"/�Z���|kydC������9����p��!�iV�g-�2u���0Ǘ�J�dba�k���TS8����p�U�$��H{Ӄ�xb�4r�%V[Buk!�0zZ�L^��fZF���D�1sk\ >Մ��7�$F�Xfl^ٟ��n�}~�x�>�3�e{f���${:�h���êoJ�.I���H�ERֽ��"0�j��\��Zk�m%D�^fj�:Y�$fF����Xp%ˈl�Qp
C�A�ܽs�s�E��8t�A��Ax��)�!���΁�3���Jz
�ͷnc0t-,��(�Ͼ��")71�	�²�è2	��Q�T���-��vk�	i��M�@I� �g�2: ���P�0���6������(>1�T�B{�Tgm͔��[!"�n�G3��E���.J��:�����Ǆ�pr �U�l�´9s4��;�\���e��s��$Z̏������kَw9#k&H�hw2 ��w$S�	䶳@