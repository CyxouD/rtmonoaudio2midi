BZh91AY&SY��[ {߀Px����߰����`_��� !������$�L�b L&����e=#�h�M��O�F�T�� dhdi� �101��&$�HE6�� ��A� 4�ѓ �`A��2`�%4��H��M��I��4f��d�G��� l��� e.�eP4T�y�?������P�����m�?�/n����1����L g����uVIfz�CǱ��pt45��Fp5qz��/8��V� ��USy\�/**�1�H�����rn*^�[#r�g��a-�t����f��Wӯ�ɄҕT���D�?��ˏgq�͛U�06�?�Z�{��U<����9�A����߶�P�89��bG��,C���	]��3�N���r񭻭7f���u;)�9�[M��8sa��
���&�ɔ�*��\��tS*�5���eg��-�͌)S��T�^��Z"
�1p���Vf�hym���˲f�pT�������j����7���j�Ɔ�䷔K��s���3x���@Sс{I;A�N��(�,� �A�)�1�ܑ-gF�u�+0�i�\vw�3�m��ڶ�"�)�kau ��ڝK�7��l���r2�!�!�T�����&g*q����lg�Z�T��3G1p�U��&��^�a�a[��O�)��ʴ0TI#0m�q`����G?LФ�k���nt��Ӧ�N���;l���f4�E[�	��;1�֘����ɴjIঽc���qt��4��-/�z�5��Efn`B	)�SY��|�~#����ꪃ	$���oZ_`�8�]�����*�KN���DEιS[!�"0�d(Bf��2e0�[E�T$ي��D�P��F���6!�CS#�����f%[�c_��|��NUU�ώ��#�ʫ�=_��??�������E��y�"���S���ۋ����$�T?0(��G��ݱ9Ѭ��]^'<�뙺B�W�|\{{C�)�<
})�rD�����^��k-�K-ȡ(��<~W+y�2G����;��cF�am?�$��R��ӮѢ\��FǤGH��qZ򴇹g���g;��JpN�d���6j��:s�/�xɔ��Ǌ!�aihdKX�8��J6^���bS����`aa(el1��ÃC/A���n!u��&k��*�P�/N�I*H��mԍ�y��F�ɂ"�S`素�5�rc���.N�NaK��L<z�L����"k�ك�b�Y�J5�a�a�{m>�A��9��p�S�cmj�&g�Dq��oS���s�z'�U��9B`��p��]�\2B1�ۋ��� XzN�p�ӄ�.25i�{���)�sn�-�YUʔU�ŵC�d����g ��m<�2#($��I-�� ��h��+�~;?�=�7�;"z
����~��0rY#(�w�EʡVyu��aS����<A<��g���;�I궳�GDjXҬ9�\a� ��e��A�lG��\.��z�a�AJxDT���lT-�Ϗ0ȣ�n� U��;wI�W
`Z��$8�4
��:B����Nc�@87�H���^�X��@�ׅL�qj(Ĥ��g�թ��$�����d����{1��H�ɒ6X;���.�p�!*#Ķ