BZh91AY&SY�"@ �_�Px����߰����`�@c�V��m@��MM���i�)�@�l����T���� � �   `LM&L�LM2100���&L�20�&�db``(�~�S��6Q�&FS�@�1���h"D���jF�h�=5�3P� hS � 7�<J g0�J�j�=G��W����q H	�X��CC����8H��*)�c�u>?��~�U����.����̼\ڙ�:1`��r��X��+�8,�,�o	^�N��d'���V�	�_j&��I"r�����r�o��Ṁ�!$g�Of=9ݏ�
~g�]8<r�Ms�b;����M�G�Uۺ��k���ʻb��v�^T(�Dt�&BM�P�E�����
�ۍ�h���)j�T^+�Ȟ��W>���[�\���Z�"k��˧���=9ֵ�4"zDYF��Ob.&�pƹi	Xou���g4��	���ՉR���F�YM�!�*o��t�u"�*�sxڅ��������ܻ�E����4*zyV ���1��A:bI�2�P\��� Q՜ʦLB5J�DPR��2J0����^d<�|���g.*L�&:�kG6\[xj�%�K�ڧ�	�-�6O'Lr�
���lr�7�����s�Ҩ�.�K�G8�g^��G�dD�_&cu޺nf4�w�/;������M=�oN#�f�\���3W�y���n]i�/�8���;��$*�fq5Y�4��F3�õ9��_a��_߇1����{d�HhP�.-u^|�k1��*��ÝVY"Ț�d�A�@�]\�.� �l�(��;�Z�_��z�ى�E;@Ё�r��S�I���͏���?YI�onz���]��|�k�7�@�������w���#������z,�	%�~�����1BI1lǗ�^R#�����xѩW�{}����(^�A	%�c�'q�#�ҮѸ5D�T�	(��-q���Ҳ�J>�'��NO�SG�tg-�/��|?�s����>Bw��_U,�\={�1�=�e�39���T�w����]M��Z��~P�Y8$Ϟ9C��E����Ԃ�TWXhFǕ��rq hڏ9a��D��<I�RY�ÎƞS�����Bp�eV��ng��n��{��CM�Nʔ����"*֭]%_[�IlRٯhDn���z\�(��-�D ���7�^���j�x�h	%��0�b��>����{y�2�^�upx�lx.�@��
�#��'�;49Ωt���$Ш����'"��M,�&�{D(|�;r�mȱ047m���>��:�t���Y�e�Qy��3K^#��l
pm�~��
���Ǭ���P��!���Ԩ~t:=n�=Y�s�>�$���좙��M�����Ϗ�ba��ty�P6�I'.�z'	���M��ߟڱJ��E@�1�;L�B �5Ƿ��Q��+���t�"���JW)�P�@�i#K/iIQ�$�p��gb���1��@��
���;-m��A�4��$J���\��2�+�k9��%z�����~��I+�dx��͊|u�|��QL�o䧟t1��ܑN$5�� 