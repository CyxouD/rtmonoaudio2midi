BZh91AY&SY�P� �߀Px����߰����P8� s��DB%(�$�d�1M�OA����2i�Q���% �� 4@  �%4�M@hh�h 4  �@"���S�#44dh� �0F��$@D�����
zG�����M�!�������K�J���P��z������&����������!�1�������=\�Go� ��t�#�������^B�Yf��e̢�R܆��CI��)�ȒG�1d�K��$0E�Z�AXʋ6P`�8P�#]\-�݈oLd�U�	B#���,{<ǿ�5�$̘�/�Xa�}x��;�o{I��A�����"�;�" 8"  �\&�I�;�X�,Fy ��A�e$���0������	�m aq�(���>gLX
R���8�G/�(Y�33]��ut�*]����0=-����ִLý�8x$Pm�Z�PL�E�OG�m
)*��G74�i���+4���)�0)5HDK5�K�[1�{���fإ��W�J[R�m��i�A�(ۅ�Yx���������R��u���� �I�I$��AM���C��Â��j{iP�F�UU$�v!�
h��� u�/�u�x,��� V�F�>�y�:@Ɂ�p�S�ݺ���S�"�/~jPǴ#�؂�@�+9 e���+�> ��gέ9\[oe�� ��]��O��,�(I1UC�����A�?�(�5��n��{N��e��IiZ2�pxɾa��S0�D��)	)��#7�r���d�Q�*\���G�:[�����Ԁ�^�j�%O�/>�s��N�2zDz����畤=�	����yy	N	ݖJO}*��[ݞd����'5�s!Dy`����+�e�����~�1	���hw��L,
շ�l�m��g��Cb�w�
�'	���8�{����/���Q����n���I=���� �>�eF�F�r�C�`���L=z����G���1kk�`>Ş[.�b�Q�K�s�#���ϧÌj�F;�;�W8+/d�Kùs�#cu�rm��"�:`���˦x8�#�X����D���lXK��2��Nl�sn�+*�yb�
-�V����DV����_�ar4J�In�$���W�!���ΰ��o�v���\�6vd3Z���#��<|˕�Y˯:'KJ�p�	�
��Gl�#�О�c���V�%`vҡp3@ݪ�@�>��a�3�6
��
S�RV>tQb��~�a���ͧ�����Z�J���6�/��ѠP�f�t��)��9�	 ��A"���>�ſ�L.^u3�en%�)�3����`���2>&�1?�Ff8��2d��;�F4r��w$S�		�%p