BZh91AY&SY9�]� T_�Px����߰����`G���8w�� I!��򧉩�<���FM)�Ѵ���S؈jR        ���a2dɑ��4�# C ��4D���G��zi 4��A�ɓ&F�L�LD��&��L��S'�=2�"h�@�M4z
6ܒA+	INHH�@�	6�r���T����������-���1�w���s5��\=Z��s��%v0����+�)x��7ʧa��L�!DA)��0a�H����j'1��?�%����"�L����&8�8Xa�b����qY�ӽh����2�^��4�=����2`n<h����ִiw�}-����$��bMw{w*�)KTO6E3]bv"��jx/����s(�ƀJ���%g���xSEi`Y%��1Y9�EJ6�K�; �%�8pIabuzI�r��S�	�IbvY��n'2�.�$9�*���6�",9�:�G2 �2�q@���o�Όf$հ�E�]-8����T3J+dZ�rʂa�[
��p�b�N��e�1naU6�^!�0������U64Q8���J�dp+"w-�Y.��3��j��N2��xm��ō���q��S��stqz��!!%ȒI Pd�Ϳ���__�Q�T�n�p�TF/�4�%)�B��8PE��@5����
���su�&Y�}���h@b�,`j��df�#5t��Vs�k����d#v��x�?|�����i���<����v����(���a��K�RMY�	�%%/^�;Lg��1,U߃�<j��C�Ix
����?�l�q���пB��H��+�B�'�3#��&Û�"�rހ�m�}�~�ې�jj.F�$S�R\}Z�`�(\�_3�����veZ�W���j�]ee�9Ѩ�힌�N��ғ$�XbB�#���|�g�Ap:`����Ƞ�R@ �b]�4��+�f�<�f1���H�oY�v������<~�G�""��<Ƀ@�RPp�)Y�ƥ�g0H6�����RD�V�PZB
βB�/�:��%��]�S3�1�cc�}'Ϙ���=t���ߊ��P��0<x�H�9�]N׽�0�|�!��И�EBZ1��#2i�J��"�;d��BB&*`�s85TA�#(�a:�9,��M��1�˨�@��@vm�k��-F \���k�¡C4)�8�q�!�֧����9��ϐl8�_\$s�D�ÏRU��<�Gbd�����/Eݵ�O_ȶ�X��uS�X�)��M(#.$�0o#��6�]-��v�#�0���W����d��Ou���}��� �2%�=���f�)ԃP�\��^l��E�H*�id>��,�WY3�z/foո�R��#f�v�|� �m��R���ɶM�q	Zi9Gv���.�p� s^��