BZh91AY&SYk7�M �_�px����߰����`�>7 �*kFh�I���ejmQ�4ma �� �� �H�F�h � hb!�& �4d40	�11�& �4d40	�10�H�M�44�!���   � DA&�y{)?%=G��~��� ���N
6낣L
N	!� �2�ڠ���
`">�@c��R��-DQBb��)Dd85ݎ[5g*|�����Ot�U���J�<�P�֘8H��_m=vA�����NƨH�-�Lq��X��yƒt����4���B"��!qyR���<7��$	�<��9�_b�&�n�h,�_��;�����a����MI�Z�0�ښ	��C!�z!Tc�,
liȈ�O2DeѓY�����,CG��-�)�ՁU�*4��� �2��#���z	�i�a�c�<�P@"���@*�����y~.��[8�d+�ɔ�����{{`��o/��6�Ŝ���7��L$�A������jj)���H�d�CC�[-i�)��s�7(E�"�Re.4��@ph�q#�Gꊻ�^f����1���By&fw2T�q��؅7����JvS냮�Cr�Ɨ�)���0Z��鹡���]M̳�>�:�K]X�d�Έ���-.�CN�Ft�m������z+e�cE�/YX̮��"$�����W�w� �I�I$�( �w�)�%/���UzVw�Y��1���G��f��BP�K���Q���b&\��Ii|�,���tw�3�"�������lI��w\h�#EUre���q����{���}�ίW�U�㿶s!�/�7�q\K�V*) Wۧϻ�Um�!1MLLYK���!ū�d	��es,j�7�$K���z�v\��C2��2�CK!��/��]�"y_�J(�J�B��h�7�!Т�Y�_ጻ�8�$�Q�K��$3�E��)����F)%�|ױ�r�%�|Y^�9�,9�o�����v�3<�!����0A��${@�iָI� ��,�������*1��(��mԙ�1~�R������UiL�Y*(��C8�Ĩ5����vi��F��\Y �B�WJ�do��m�AA�t��O�4�Arf�Ĭ������ŭ�5�y4�J3]N�$
������^��`?
�9�q�8x3�:�\�4���ǅ�>I��0�ؚI8TF�uE�h5+�P�CLh����v'J�ҫ�Q"(.b�8}Ўʤg
��"��*�A6Q,��K !B�G�� ��n$�`����z�-�>����H�"k�vғ�H��l�k�f�H�����h!Pb�[(��&���Y��2P��i΍��Q�sT�%X{b�����h���h�9�:��t)ċ��í��RVMFJ�l)�19��t�(�H+��e�Bd�k'�8�g��m�4��i���I���G�O!�\���Ӽ<�}��S96`Ob�E�ː�c�B�2;L�1���f5���2F�;���]��BA���4