BZh91AY&SY�� _�Px����߰����P�8�@�;m�M�n�$QOS&�i�i�<�=&�m@ѣi2bO@ � yF@ hdi�h �$��Ԛ�D�h�  sFLL LFi�#ɀF	��j��	?F��?H�4h��244h�G�@�fK$ ���H\(������B8vҨeLR�����M��$	L`�X�:CH��msr-;�O*B9�X�rY����هM)�s��A�TܳVaX��I���	&t���7����)IRPf��68��Ye���d�թNw|�6^�!Z�(@�1{&���o�Zilq�{�^㟔�νc%:[,�v���!�I�a�Ī��qNL��	j/W/�m$�yX�&8  ���P�	�tWH�w�j�h1�1YjF]�;q8�)$��7L�Ŝ"@$h#�Er K+��m��I%"�	v��������튒���+W��Y� ���4��6�*�� YuFr�yLDH�PH7{�QM�R`B(`��seʵH���g�����xGP�	�Cm���DM�{
|����rU^��(�2Y�#�5!x���ndV�@UQ�$��"�b�b�aSdԂ�alat��X��HDڛ���M4u��U]<8��>K��v�1�߷>�Xӗ�֪
��Ն'5�W��R��N?xd	��8/\.��%�����d�U��t?�e���#J��oHt��CiЊ�������s��;��^�N�,�|�$�!rvG�]�Vn5�3.�����S�/�l͞����(ژl�E8
��vl�c`QUk����*䣗-UQ9-��p���:M*�!ے�6tR��	d�01k���N�Ě�;�Xu#���l*5V��!β�\�3ȿ���l��]"SxJ���R�I6$"�VkZmD0we�"`�"e@wa�t��6�V��
v�9p�����ixɌw-��F`y�=�7�8l�fQ!�661�����D#{�T��c4�5[�F!,��s/8B8�$�+��H&<A�ED47�#��M��ƌI�N��`%j}7̑�0�8tB;5H�XTWqU7��&�%�Gu�,D*�p�\��8��F$�eHF�R���+�7'� ��zS0��u��	�d �Y�H�r,}�H�E�C��*bƐ�l�9"�-z��v�"��=(7yۂf���Η��Mh
��c�Ė@��C�ude�/=� g�ZMi�ۋ\d-Dj�n�P0 x��RB,i��D���r.d** �r)W]���}�z�������)�R5g��1�4�Bꛄ.���R�~s ;$	F��2�P�w�-����4�7�l�*���"�(HPm 