BZh91AY&SYA_%` b߀Px����߰����`O��p��%R��W����M����B'���F�(� �(   4   ��(�  i�     �~��2 0F���@ `�1 �&	�!��L�����D�'�a�I�OG�2�@m52h�H*ߙ$�,$A$	9!"��o��` ��~�*2�|�@�0�_R>4��1�w0��V�սk���0uJݺĳ�
:sr����(�iV����'���h�	$�l9A��l@�>0H&uF�H�:g�|�,0�F;�L��&UWM��a�RW	�]��뻽����00x�xSu��ϕvJg��f�[vt8��fx�΂Kd�K��sl�.�P��iZ�^��Rm�I�P���.2�V��Zv�(JP�vv,h�vÛC
֎�X�C[9ڡ��K ]��V�T�R�FY�N��+�aFNB8�dg�Ɉ����L��#�3�2�j��X҅.�SHVDf����!Ļ�\��ю2�م�(G�J�*r16�N�dJ��1 �U-�U8�!Y��ڋR�glw1Tf��n6�X(.j�ٶ���,�{E)gT�%�!p��N�SҘ�k�6.���5��D=� �)I����?ƿPh	 �I�I$�
@$�s2Q�WTZ�]3a�i���LQ����`�C��R��tKd���CH�"� iw0�gk���Y������Z�3I�
��+l[��(�%i��O����8�,� U�����}���Xz��щ�,*�G�H0l�<>�Xq�@̬I�
x\W�w�����Jۏ�{�}�N�g*k^���g��B������<�����MY��ǩd�%6�;�C#�s\��4lі�����_<=� ��/��CKQr9�"����u�)H{��]��s������^��Z`Մ�_�4�P�w]53��4$y�,��$�� ӥo�*AM�\�����̩X  o���PG��c؂��#Wl�zf�ROM
u�� �����\��B"�~���A2�:a�ʟ$_=�{w�	�贛������.�x��N"Y:ʜ�4=��m	�q[Ϫ�N@ˍ��z��� n��>���S/[N\�'FVI��k�P���'c��@�} ��k$V��<M��I
'q7�!&��DPT�Jp�tU#^���*�Q�2M�%�ݗ��@�B7zl	�ᙩ�A��"��>2�C<*�0yuyJ���Ϲ�pAY���5p�6J���!��u�%ic��zT��i�A��4���~$���5��JƖA��N le�6��R�j�ݧ55W���}��J�	�`��)8����	����2�ي�4�؃@�\����U�R�GJC�)83�H����K�V��@�A��rL��(�9�3fpo��#�j�,K�������H��;{Y�2���ܑN$W�X 