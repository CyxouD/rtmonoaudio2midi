BZh91AY&SY��� Y߀Px����߰����P��4M�ld��!$�d�S�)�Df��=M�=OQ�C4���?@	J b� hh   HE4ESOPi��2  � �����&L�20�&�db``$�L�OP��Q��҆��ښ h$-|]P�,@"@IA'�{�*r~8V��6��Q��.@㴒U"�mCH�Z�Ȳۻ]��%��S?0�n�w��OLv�Vt�%�]vʡ��%�*�tH�]�[*�u��g&��nkVHei�q��V�He��09�_z�қ`��%J]$�EE����=g���	�Ɵv��x��O���h�[���A��.O1�ȁ�9�,)��'af`/_�yH ��"m"�.0VC��AP�V*���9��(��B�٠B�Z�f�e��R*�*�[1l���l.�Z-'jEt��N2۹� �ӵ��`�j�(�V(*�2�-,���Ħ)���jDHl��Gaj�:[��*ˤZ+Z�gcnM ܨ��r�:�U�T
�0��k�/2	���W��;$�H$��m�@�
ǋyW���^~�K;ʸ$�)�2e�|�jbZp���&�Se|��b�&���(�4��&����3nB��a����{.F�a�[5���]��U]Yaw1޺e��va	�x������N�?*���)��.+�S��y[����*����N[L
<�#�����xѬ��u]���2�cA�a+:îM���P���s0�]�kvםcr ��ʇ��.O�tIAѕ���_a��@}g܀R����˒Ѣ\��F�H��z��e������)�;��I�Y<�x�����P��3�p`F�A����5I� i�wH��Y�
�Q�����8$r��)��f���1����$��*R�*+o:\O�4gvH�t��1��D�jG
2Te����!��=-��ӷJ�HAa�D�b����>ŲY_���x��0׽��n }"Wt�:����`.8X x�ƶ�#���<�C�"�����h7��l��o1�:&���Z��PMW�=������3�#��F�h�f�K9J��)�\�Y@ NQo�&��az0@,�wA$t��P�
�D>��~�S`u�r�;�3`�6�f�ָ:�#��$dz4��m�hat�ߩ�0�p�\�x6��4>����ʌ2��īV�`3E'݅�"�3Zw��_�&�^s���%=�%c�E).�aAQA��Z�� l��vT��sO��ѠP�����MM���xI'	X6w��\9����S9�eڒ�MR�gy���2<L�d��8�=���3��4a��_���)��(58