BZh91AY&SYc�(: 2߀Px���������P��Ʀmf����I CHѥ6��$fP6�A�421�D� ���@h  "$ȩ�Tg��i�=	��@ 4�0L@0	�h�h`ba"Bh$��=&�#i���#@2���@���!
�$MA �P$�N��Gww��UFZ��E�Hj}�N ]���X����E�-kf+ͷ~В4�SMI3�������f�)VJ �"�d��8�8D�H�L�2�@�l�n�ѩ�;�uZ�#.2Ɏ:\,0�F<H1'3Xֳ���g(��1n�h�ϑ��Ja$3�n��w)�q9������-��g�s7j�"Y�Q����!4��T���NC�{�@&�&�&�i��%2�aqɵ�	K0�d�vQS��X�+��y�Րp��¦y7p�,�@����4������<�eH3l�V����k&�֝�Qb�$FbS	\�A8�V"��;c:db�F�^��}���ٱ�������J�`PI��eO����(����m��4� �k��������r�J�i�"̖qX��PP},0�%�ʑ�h����%��X�XI\�*c�Gl�jaT�֩�b̘�m ��33Ǫ9������ˎ�8Ϛ�A�ۂ�S����G���'o�Ɠ	{�U�6a/z�ΩG]�|���ل19�/�]�#�W���5��m�_A��ޒ�1rI������n���QPjhlI n'�O���-3E��VhSH[NJ�:���J��c̀�\���E]�A��Ɓ�QTpJE��ɫ.����Z�^�G7�J�(�ckL౿Y��u]��4���oی�H[�)jX\4 �#X��t�'�PX��aq��PiQ�	!�̶�3�W�δt��1�ê�zf�L��RP^�$TG�2���;,���L�Dʀ�!��z8k�W_\(>=
r�����l�b�L~!���D�1}�FX��Q�l8A$Glc�O|�n���]/���f�[K�ZD���\�c�f��7��0�z��!��t�/�\OXi��3(�I��%j}��HD�eT��g\#��
�5WU�("a�Q&hu\�I�����\Y�Q�G�4r �u����W�!�����i��I�0o�����ش4���p�|ح����!I����Pa�IQ��sy]zf��,�b�`�g� ��iѴN���y��n�gB��7���5c`j�۩���0@�{�z�H��"�M!�����؃!Ъ�=W���{ȋm$Q4�3,@�,�V�f��\�g ϶̥*Mm7��Lٜ0I"��E��2���ٲ!#�����6�f�j����"�(H1� 