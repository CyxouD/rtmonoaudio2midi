BZh91AY&SY8K� a_�Py����������`zI��;��Z %D�=OQ��g�4��@�hIP b  4ѓ@  dɓ��&	�F�!�Jd"�4h  �  �F�2d�b`ɂd ф``$CD��&L�����L�=jhi�А_�ܒAc&��!"�|�������|O������J2� � @(h8����LHE�V����EL(�g����A�%ǎ�L��ρ��.g'[V��쒗��j�%ZU,�9���N���"�K��U���M���;���N��樢Di���'Ĝd�	����,,�?z���!ez$$%���B��9���zR����a���.ݻ�}�C�[}dVN�{��*=�|[��5�q��1�;�Z��2Sg/�I5��L�+����,H�ƍ�*a�깻�i�$guB���tJ�DmA�F�ki��To`PH@"J�6x�q:�	j���TN�!���-/
S͛K�k���R-�.�'�HRp�P�(8U}X�Q�p���vS0���Z}���a�S�A. 0T��Aթ�,�E�2����CА�zp-�eX�e�4>H5q�o3l�"l�ۉ
�-v��G.�SB��u�h�PTN%f�o:�j@W1nQň��&��+��$Z�x�{��8A		.rI$�@@1��R'�LG�ѥ�j�y�"Q������BJ��2��@_ɗ���S)Qm��6����V��0�Ux�; m!L�^��G},�)d��m�F#2c���Kc���m>�͒ߞ����PM�->��'�-��;�G�D�� ea4�K�D8�����!�K��#�q�P��jVz���>�.�P846B7��'y��[���ȭ*��6�'	�c ��ܼ����@2]�	3�iSg.Q�fj,F�$U�R]Xe�)�����S����T����R�_Mf��,��N������|�`#��Q(�B ;�$*�Rl�W]�U��-9o**��B�yS2�Y�e^0����M�.+��Z�����ҬzV����unҘ4%%�A�J��^��,װ*^�}ք��y@]�9KMzG5�Ĩ���7L��5��Ք� ����ǌ������%o�MWS���,���HG(<:�ha_E�[���\> �E�4�&�%��ə�1��#14�%sBj^�30QE$���o�#Y��)�Nf�RL�'��1�0@@5PG7u���7��86 �Qb��̢�4�k�Z����͔j�Z�ŹPd�C
V��D#�t��d��$R[n�t�I��9�0=� �ƾ�'a��نC���W,R��Y��2`A�9��0o�)��6U�V����󚲜*�BT��Ջ�{���-��XX+�bf++o�"��� �9��q�����J ��&�]�ۈUz��L�<W��5ᴯb�#^cn�t� �m�Z��S�d�8�$li�n���B��]��B@�,�