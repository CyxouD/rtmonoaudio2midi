BZh91AY&SY�:}w f_�Px����߰����`_z�s���D��$B�I��)�S'���S�M'��<�����h�Pjm J�`       "����L�&�1&�A�4!����@� =G� h  =M � �`�2��H�M	�!�&M�bz�h 	� }[��&!	@$�O�{g���~S�q���C ���~&���ch��EY�=k{�N@����e��8z;AqgZ��)9	)�d���&6Q�R-���UtU�;+�C)�dKI�*�>m�2
99@L�$��E�]vzO��@��a����wgq�x�P��M6�m�~<�ŗ��N�Ǡ���	4��ե�ڃ��3M���Bͱ�y�8�4F�-��Y�������R.����q2�S*�2���sI��[M	��4���(�5�G"VD�,�yo��˭նٶ�$3K�oa���0k6�y�x$�Pl�àH8U �	H� 3	Hl��V�٪�#P����Yj�֧!C�&J�5�4�.]��e���^����$�������BKp�yM�,b+����T�!*��u���n�(��"������s-��ˀ�ӫ^���33�T�ܹ~��ϋ�mTQ_����E�{�_ry��q����-7Uc��$3]4R�JM-�}�1~)�&���@dk�c��(W��af���� M�,q�C���h3�ӁD�	,g��T�@���蘺�[`�:�2&`
�e[U �����W�H�ܭ�U7�b\2��ȀҬ��q��k��BKN6���6�R�����`@�J���H�7==�g&IN��#�ռ�#�S����1�j�}��@����~��#C'�1�D������A�^Z�߿�J�O����,��Z(ӎ�����oc�n0�$�a�A`Hs��a8'�
���/:�)$��%v�L���kk̃1���D�zL
�z����AyM���.�;�?L�ݭ00��p� �Th��`�a�$7�]�(%��vaɉ��#��#�[X{7D��D�W��S�|#�����g�����+U��0	�Aǂ��F�7�:�&��a����.!��$+��KKlcEdFDө+1!&��vD�LP��p�pQ"�YM;�(��("a��L�w/!PBR��0M�}��ҁ�7uA�-%Q��A���Jú�^�Y��-����Q�9GI�r�f�i��@�1�B-Ġ��k�@� �NJʧOav�X����jK�ʚA��I���a�H�<y���*�(�f�Z~�S�2F$�KhW,�~��Ċ������D�ڍ��!J��2�<��n�t�X�\��)���V-��MQ�;�ǅ�Iܨ�tay�k��D ��)�O�V�3�2F6?_[B���]��BCp���