BZh91AY&SYj�� _�Px����߰����P�8�F\��D�dИ&i25'��Tz4d�&�S����aRhL�2dh �DF��   �   9�&& &#4���d�#R�MS�C!�M4��444ѣOQ�Ԩ�>�`R�PU�����Y���&Ϭ���IQ!�簵(:��@$����&��4��{���N*��"Q�ߙ%n�뜱)7i�3�j{)Y�t�eQ4S�UU9s2*�l�����QD����	�Ӎ4d��cxen5���w�7���3T�n!�>~c^���D_f:4r��KUXCщ�m@��6v;����6BC��ԏ�tG]y��4ۻ����ڣnTP�de�3ե�1������EE�g��v���#,�p�2R�����'2Ʃ��5���=s��<%B(�Sy�<M�ʳõ�!h֓��#S6�eb�eiH2# p�����J�ErjÈ����E���%\�� ����I�`�R�.uI&�Һ	��k�j�$$��$�7�p������2�OwD���Z?j!Fh�ܴ1�B�DCR!��ҩ��@��;��[�a��G�^� �X�1k_��3��NU�۟&,r�#��^:'��1o����uh�}>�L�g�^8�-�*�B<�l���b�W�C�B�)��G�ގq ;���-u�;=��2�c@$eY5���o�~G]��cd3$#�tνy��87�_Z͍J��!��.'d��>�L�ݫj��i����!�K�c]�P\��GL#�P]�[ZEf�������N��픡
���]�#��d�j}�^�	��$0� L����kg&���2�ZA�`�عg�4,)ɟcd���H11M�=�y�8�2���Q6���a���k�N��vJՠx���k��ɜ����[��U϶\6���FQ�Y9�:F.c�7l�����N#@���+�|i����W.�}�l�bp��a	kHG-�+��ۅ���h:(F��$; �&�(�B��
�怈d(�N[��A�`�f(s�|���8E35¶h<�R�fi.E $:�>��6��Kё!���$�2�FY�!������f�A����`ಲFa��o;6�(0�m5�oLA�����RBSƘR{|�I��aݣtlY�8�^a� q�́DA�k�~�]�<&�f��yP�<"*�F6�WU�H�I��6y$"�HE6�CE>z�Q��P���PR�b�u�c<c�ʆ P<%���2�c��x��n�ճ��v������8y�	�#�gQ����c{�F�L��h������)�W���