BZh91AY&SY%� $_�Px����߰����`?`(P
	$I�����&���yF����4�`j=5T��%S� 4�� �  4d���`F�b0L�a�101��&sFLL LFi�#ɀF		�d=�$ɑ<��h�&����A���	��A$� $\y���_�_����0`�"�@5?o�H�|�#!�,����E�]��ˏ�fZ!�S�,��@]��tי��"Ң��i���6V�6�Ү�HsRh��	h�p�i�sA��ӝ�lj�����q�p��	� �N�Y�����.@@am��%�_A�m=fܱL�00Y�Y2s�2�豶�"ϼ������S��z�Тke\	L+��҉c)[��IvR�*S�X� 6��@��,-�S�C��-\��[rj�,#�:w*o�i�qUvrk�r�ʾ˼f]������+�F�rRQ�$������2�g
��p�9)�鲹��U�;�eT\�k��6aE���v�IG�[EPi^��!�!�Q�d@p:�)kH\+ v��FZ�e�*�n�~]0��YBM���	�#,��:��$�N��S
X:�E�6C<0u����*_��}����m���ɶ�`Ā�	��
~��?UV,�tF�w�L�|�"���"�D��%X?YH%���@1x�T�FB����W�������*b�_���QJ\�.	�~��k|2l��yz��_�y%e]ҭ�h���QBd����Jw�@1�D�|�W���Τ���R������g@������<��A�!x#���27��&�}[���h���I���|�x#�:�+���^��@y�P����c��h�YR�����U3�4��>+���y��^�;s�	�Vw�4��c�Ij�l?
�gƐ1C!�t�)���k���:�:��#�2�J�J��1;�4ZP|�]�\��Y"�]T��T 1+���#��P������H
Q@\��T�v�V��߼���Rߨ�/g7Q���:-��P��=\hNkf��Y�!]\�lc�/��������_Ŝ^��C������x���̏k��@�}`�4	FT'`�-$hQ;v D	���Б�.�8~����b+�,UNEHA6Q,��^����V	��.	���ڍ�@oB��3ۀ�����������8��R�AQ~!����Z�i�#�v��[�F4 N��Gbd�g�6���
�����Ny���lKPw]i�,�T"ނ��7�����m��݆���j,/Ƣ��Mk�����0$��=��šl�)T�䪍l�8h:Z��!�~9>�/rC !.���}@���_aC��WL����O���O�I���Yc�]@M�j����[;�T�pi�ȑ���.�p� 8K"