BZh91AY&SY۩0� �߀Px����߰����`?M��*�DJ�I	�6�Mh��)�S�m#FCL�4�jm JT`       挘� ���F	� �bD�� �� ��  hɉ�	���0 �`�0�" ��S&4�@F��b4��h4���ԑ 2�n��A�$R%���� _����Y C>�~I �`�1�w0��V5�Һ��2� �ۦ� /�
tǶ^5�0hK0˪��`53@��n�j��K!��Z\���]���T$f�kю<\,��F63�=�8��__r�\� �v�I1~=��g��&@00e��Oe�&�Ҳ��i(Ao'zmѴN�;2�X%���,,4���sj--
�5%�t�:���2bBBn( �è��?�ί�[ܫ��<,��w��t�m���B�\}�)�&��:p	��ak�[dT�Kq��H{�h*�	5�#B]�]kFcN�^�^Ӧq/��9*˽̘���L�2њP�ЌPia2�,� ܨ�[��P����Mi,��::�P���H�"��sYEW�M����(��)�M���C"k�j"��[����=?��r"'$�@" w�a�#���&��U!��[c�a�B�݈��4?ݤYQ�$D�"a�gH� 1w4T��E��2��������b����pQ�>��S�඼���T���G��������d�)#����M�/i�Պ ?M���~3Vڈ�dN�з��{z>�z�:Č�,���?s�^f1��e�!���a�z �@���{D�:�ʼ݋�b,�}�$��ʝ����tϿѓ:�Ǖ���� �K�9u��Ƣ��JF�S��US^��Q�0��^��G��%�ug{��Èӳf�iV�ݴ���@�!�+�@r4���N��MT��XrGQ�˙R�"P �Qn-i��/�5��e���Ħ��eE����z�6�z$���������PP�9�{q�q�
]d��%\Hه)tǄiV$�Q�͈4[)%
��jLb &���1���a�]�iὋZ*��& E� �n����"mkZG"�����P�m%��;F��i#B�؜�Sﾄ��������F"�Q]�T�hK�d �(�y�׬� '��&o�6=4# +@����a)���y�׏�"�;
��A�9�UӘfK$p��Y�{w�yc@�ˤҙ.����U�o��/2/D��dӪ��k��0ĠA��o+@�z�cu6W�0ջ�Ί�o��5Z欺)�.rK���] � [=*�[��U�
nA��Yk׫Co9>20����AD�f>=�y,�?QC��W�' ���[Es�x�8��������q�ݘ���%JF�"�n�'���"�(HmԘM�