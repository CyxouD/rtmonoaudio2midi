BZh91AY&SY� �_�Px���������`{w=�]��❚��I22�Л*y��?E<��{T�hi4�CPj��U20 &�0�	�&&��Q�Q� h�3Ba4� i���Jm� # �2h�L�&`�1 �&	�!��L�������F�S�$��螧�4�L���2	I e��H��B�$	?#�_! ��.��G�@P���"�@f6���,���.^�L�� �*��K?� (�c����ܻ�H:N��Q��io��H�q2L��(��D��2Z�Њ
%C"��Q�<Hf����[f ��
�T#gN�cE�v �*��j�HFB��9���ym�a ����^v{׮0��ܭՐ��Ymkm2W�DI_��m_}�ݙBCl�ᑹ����� ]/U\J�à�1y��*�A��+�Ȏ
�^���W�y�"�܍�0D�$HD�� ��H^�r]9�7f,V�f�u�EY�\ښ�jFQ�(��̦�P����(M4�iKwfH��x�Ⱘ�@�u��%�4$]2b���x�v��3ՠ��%�6�-\3"��\`�Xvb���i������krKd�[]f3�&k4�!0x䖉2e�����ot�I�qp�셴�&���8Ħ���!�����k��홋��	ި�B!�^m����A�	��t����Xն�m	CSM�;(M�	�I����uR6���ky�Mf�b�<�E�.5ք��qqS����ͤbsl�SS�y]1�Z�Y��ӌxb�u<YOĿ�<P�nET
��UL���^�527'1)9AQw�#of�d�f�����A#o��m�i A6�}
}�����W)`�8D]�λ�7��_&�ld��DA:ؠaFA�K�KD�� 4�l.�A�tw�`�{ML�ěI	f��k]�w�5q#Uu�i�=�Z�j��3���yg����,>_>�I��xJ�̳|��� ��χг.d�	8�����W¢��ߎ�Kh_�s��W���� 9��n���C�!v� ��؀Xl�q��plx,�CҏM��B�I�H�Lr��b�_���p�
���c� �&��#]	�
�Ì��j���7��ŠR��^��V�;j�-��g�F�!ۍ53�Fىb�bH�#�:W	2����=&'���J�H�9��br*�&�h&0�VPu	�)YMrT���X�J�A�p�gƄu_g7�0i *�+j|Q���7�j�y�*�� �oщY�{���X�3K�O5	ҵ_g����@s�cc�{Oրn��]��8���Sh�-��A�@ٱu��5�6�N���s�f>�uE�h5�+�P�cLh���(�����&��DPT�Jp��s�#`���*���e�n봰�
���{�:H� � o���>��ߧ��&�.έzK������9�Y#@�v��Fɰ��@۟B�2\��5� ~�M�gīk2�c
�T�h����Iõ�|��i����ċ�G!�z�8�L�X:���9*Z�J
Mr�Ԉ � ���қMj�TT8�3�T�ddi�mx�Ġ*I��zE6�}�y�V����8��A�D�MEIȾ�V��� [G��V���׺[8D$ni�o�u_���)���Th