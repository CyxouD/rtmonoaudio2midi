BZh91AY&SY��� _�Px����߰����`	�}o���D PP[�5$�	$&A4�F�=5b��0G�ɓ�jS�"�I�4�� � C@�4d���`F�b0L�`���44 Ѡ �4�Ѡ"�S�(h��z�4��2h �F�$��j�#���b�~�zFC���Ad ^U �L U �P<��&X�AU��Y�
 "(V��?�%�D�$NP*)x������I%��ϧp�?�48oh�i��g�OǺ��{׋��Q�HaչT(�썠�E[�T�ې���j��7���1IH�l�)R[R�������ȴ�gN��YDT��$Qd�RuI�iJ����b*�	Tꪜ�-FW��E乙�����_f0��Yʔp��<�l
��|��м�YUC+갈�����U�}���,���iUV���d���%��(�����8���ٓ���,�&�4\ܭ�Ҳ�Eӎ2��ZY@I�WqZ�w�?8���U�޸yn�O]���A���H̼��{`57*�e�Ѡ�՛Ƈ������O�s^����;;�d,T���-!b΍�SO�'�p�ctԧ�p�oT�Yg[�Y����b��6�0,	��-e��E���h�6؜j��ل�%�>fhյc1fJf+��p�q&AYט�����}\�-M\Q�Q��Y��}*� b�N���.
��3�ѽs<��&1�Yx�ޞE�n(&b�v�����U��MD>�U���r�"{ٽ�߄�2+�KZ�'(Zb��f]GW"�9��*S>�Lʳ����Y�2:$O#��D]�qvf�s��7�]�e�ʻ�-�P$A9�\�9N�U�r^U�r!(��	1�� �ed�Z8��U����.�������v���QZ���՗��r���r�B��yt�)�3��5ɱJ�s��nq⚚5��0^q;*��)t`�9]閲2扮��Dt�u�ʰk�HM�ad�4!h��j����:��Wc�էk���ij�Foh��]@�yh��́@*'*gnܧb�;K��U"���7Ғ#�N�i��;a�wh�4D\M]fȔ�ý��g�O
4|���
��ٝoȹ+̙+-���k����0uP�b��s%Rw;F��)֛ɮ��I�9���ܪN�][�x..=�yG�$�}�+;�^�4�Ni�1% f-W1��v���QI�]�z��6��975)#F΀��C����oM����Q3��̧�&��SZi�f���=ns=k�3�qw��kJ�|Y���g6�'��}老�� ���ci���L؉�.9�4'���Z	��)O:�@�h��4j��KT)IE q*H� z�E�?�R��� U`�se�-�끓8��;�LVDu�p�7�W)��NT��<��=��W�����O��o�/([��������w�MO=2.�o0I%�_���L5!$����g��=~o�#ƍJ�p�3�}$v��7!$������M�rO*R�"U�I�9��W/Gū�	:��e15�;.���Jz,\���A�]���%/�X��^��#{�#����u���.����s�.�)�;�t��ڮ�AT�d�l��r�.���߅N-��Eu`��6��C���Ds-=D^	$���m�Cv�]��؆���'1����?��
��;���}��r��EV�h=%���r�5f{�vl!�=-�&�-�zƅ����������Z��Q��I(��Sۉ��	݉Vӿ�Y�C��ck�vl8E ��������۴힉jLY:�b���0L�ݹ�9D��s3"ڢm�1a0��e?
OF*h9�9JŶV���Z�Z�'����8�uwd��l7��	$�I.]d�vi����
�ywyN�����;[d5ɾ�p�����E9�Oi�v�\�
�Ꭿ�X'��2���7��N=���v�[o�۳�,R�uMba� ��r�B �5�Á�1��͂�N����L�*:vYr��j��BF�:m�<�U��}��g�Grn�6Ȣ�X�³�5gmh��xH"	\6�EX_4�˙\5/u�8ߡe�JnFx�h���I\3#�f�&'��sٍ�w�#FL��vj
��H�
�C�