BZh91AY&SY��L V߀Px����߰����`_-�� �LH��bI����)��oQ4z�Q��4yG������R        � �`�2��i�4�h�=&OD =M2 �@9�#� �&���0F&$ M&����16��4P =F5.��ʒAS&��!"ā��S�_ {~TReL|@@�0��$��1!SGsi0�����{� ������)ᦖ·���g~�3��6>�vnD�$%ŕ9f�*֋72Sn��B��ʩ����A=T�H�(Y�spC��4hjP�cA�.���4�?rB�7$�R�BBX�p瓯���*`3~<���gV�|ѿţh4���-]�he���]Zl�f�����qj��&�K'���+臌'��h�,�$FӇ���Y���dE�$\�/���+5��+� A��� `QE�@�	O�u�v[���d���5F�i�sMÍ�mB�,:a��0e��q��Q�0^6��R��V@U,�U�ˌ'T����fb��!^�G��7AIA�QjABM[<�[T�x�c��%�%d8,Qp�+�1a�R���**дLGe l@��"1�� i��J!��]�����17��[�J���ZV\d�f��qa��ꭞ:����ƺ� @x� H��&���;Q;T�q��Z2�N��)v�@B��,4���J���I���D�%qDT�XA��ך�+X�;̙s�P�bl}���y,'����WA�XC�}o��l(����m��w�!I�F��y
=3\��r��p'�8���"M���~�я:
,�_Fð��b�b�4�M���o�bp������l��M�����VV�қbs���WI�<�G
��h\�-ʀ��Z��ے�1�=cFcd�#C�#�R\p�+�(Z�^��G��%d�u�]r��������ϒs�P�Wl�gt�h��2M D���:Y"��>x*K��Zv`Pj�) ���X�ci_�0�Uwߦ$��\Uu��5���2�ܢ�/��e{�&	I@i�(�F�-R[��L��������P]Vg&,9f��7���F���g�fT�� AK��ǔ����J�.�]g{:N���P��HG0<�WpB53�����\>ptEd4	
����4Ɗ�Fbi�JƄ"Ծ��0B�$���D�Eb�u�QJ�MA%R�3C�x�B�F�
�=]X#@5 �waZv�"�������xyXo��a4D=�us�J��i!'Aٻ+&��� ���8? ��B�]R���⽘\}ӵb���Z����PFܴ��F�<O�i�z)o<R�.���5�q��[�u�{�X�ξ�X�AK����r�1d)VA�s*X�}��Z���"�	i@n&�Vג^���3�y���3t�y
��g"�e��6ā,��Z����\�cK��s&H͈v1���_�w$S�	����