BZh91AY&SY��0� _�Px����߰����`���( �$"TJ�HFA4�!�F!# 2dh�5O�)R        ���a2dɑ��4�# C ��j�DMMz@2=h�F����a2dɑ��4�# C �!4�$F�Ҟ����&��M��ɦ�������q$X�0@�@���� ���{����6�$ �0��M��MA��1�pa"�/k͹]ц��@O\:b=�'44^�ciN���n8�d�N��a	#q�#wm����E%�D�9i���##�jۤ��Z�v���[k�� ����&��8��+Z	����c��k.2ur�O5B)E!�~^��\�$����O�7�οګ٣+�8eu�t���Jw�<�%�`"A2�} �B�q�&�>ϩ6"����W�e�Y�UE�'wR� ����&4i�+gX�
�7U�"�+�̅,��L��V@$Ⱥ�1g�y�IfOL��p���+��.�v����e�2�H���
"�x�zS�e��.�Т�8.l�ln@�<���S#.�)�=e�Ƙ�B���ؽ�W9(p56	�a#�S���Ɍ24Gg�&��t�(
���!tgN$���z+3����Њ��:�=X�E2NԨ��Ni��b�h<$��]p�#k������0�Ιd�I��U�q_n��^T��w�d�;q.;�s�GbA� �j�y�H�=�9�7����wn���p�����sV+i�1�o{̈A��&�P�X��ʐV߂9��s�93X��h�|7���'k�\1s�н��Z!f0Ayh:[E��Y��R�6!�;�Ҟ]W��U�N[c����ȵ �� BJ�M5x�w*�����o�Y̯}�
��ތf�t�EU`It		M��l� ���e�D��H�Q4�������,�U0��z�X���3	L�j���v�=d�M<�n�x�[�u�p�	g�W��������9a����ۄ�];�I �8>�����h�Fv�wm�:|��t$:bc%�ρ�S�p�E���N������H�nhm$����wH��co�X�D�Z��!��"���B=O,:�ҿ�� ?��I Gޗ��N��5�z�Ղ��{�I.�l�t�J	��^��d0q�F��r�;����8`@�{ި$D�	Nt��g�Ap:`�9c�A�4�� rĻñ3K�.O`����H�oa�vW)���I X��6�Ѭ�&G���Ƀ ��G�e	#�|�|��ې�4��ad��옴�4(L]�Nh��������M��$�)��61�I����4"V��L/��v䙱�ŵ��HA�$�zڹ@��gb���τL1�tEHh9I"�S%���t�Кw��@��¹�0B�$���D�
�4�EX��&J�g#��. @9L��&ϲ��\� ʒ ��E&��P�\�����A�#O[�*����9��f��JL��B=��n�W͍$ �X�B7�I��7�פ���;�:��]&\�ԭJ��Y5���kə:k@����sώ��{���욭�h&�bE)~J�K+���Eƶ��U$f� �,�o�Dh�R�c�r�Lo�qs[�:R���D����=�kN�(ZY�7�,�F�%C���F�| @`fG�̦��ŝ������$o��_�w$S�	}�	p