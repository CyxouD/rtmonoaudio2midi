BZh91AY&SYT��� �_�Px����߰����`�[��j��%(H#@	�D2Sz��L���I�i���=���A��Ʉ4�M!� 9�14L�2da0M4����%2�S2�� @    �A�ɓ&F�L�LDA&��==&M�L�� ƀ%	/WI
�H�HBBK�(}��~ B����Te�6����0�ܤ@�h$%��ch�a"�0k�Z����H\R��rY���;���(vj`��;�|\�Kw�XHD��	�'�$!TfZ��kGJ®�R�W�D�� �[��v���&``�e�N8�=�����mi6�v�9�sw.����}�4A���z�d�+k��NCN5��M�7�-D���9tȦ�)�UU��U��f����	� ��
Xa����Єؗq�C �ä�2�S�	%�2��������EDMb��+�J0I�Bb�
�*�)���uӲ*�N�nWMP�y���2�ic�ۨ���F[%y3bZ�y�ŵӡ����2�?/#��r#�!jԒ� �6�α"4tKM��Y�M�#���dز�v)�U�Lލ����`�X��T�eN�-�D��&Z]��ա'gI���&�"�"�ݳ���y�Aڰ�)���K���*�Uu�t2`g&ݣ_h����~�N�E��b.��JPxXʃ�3ڨz�Ɇ�D���7qi���m�(�l�z���L	!!%ΒI PC6��S�D���sU\���戻%��7��Т� ����4��l�����PA~b�!4��Z �tw�`��[7����S1[_�w���%=4���oI�vO��KO�
�=}��я���1i����u�W����B�g���Sn��($Ӎ{,W����RG\��qe�yO}Ν0�P!fXeg�;y����RfC0_�fr��Vt�]+5��R�)����Ϊ�4���b�h����S�Kя���k'N���"z��[R�3$�,�^<��ww	J	۫�w���Y�:��^����v�S[=4���.Z�i$D��N��L�6�`u����TiU�	�e��&jĿA�^$�2���%7�d[,T���*��"����>��� B{Ӄh�����6�6�!��!�I�ag��f|��B��I��-nP���+���h B�W0�0׽��@n�8�2�1�ei���[i��K$���B�ع�PЎj�t=�a�����"�	�cE��E�84!(S辒DPT�Jp�B6�#`���*���e��u�, B�P�N��|��`p��������P�[b�?�T�9��W��͍�Z�`ܤ����m7쵅(0�!=��B9S%��6��{ B�^��Ǔ�_�.��U�T�����1�;,+!vQ5��F0�4k$�^2��৖���C�V�VЦk�	,p��,U�AM���UF�B��,��j�~z)m�!�:N�&�m��[9��xxR�A�}���RT9/5jp|��
�dygb_<�^�ms�4�d�u��~W�.�p� �?��