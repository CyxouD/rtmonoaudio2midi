BZh91AY&SY�1$  _�Px����߰����`o�ƀ!��T(����BS�5'�D�'�d�M�26��� �� b4 �� `LM&L�LM2100���&L�20�&�db``9�14L�2da0M4����$D�2jm�OD�Й=@i�$H�̒H���$����	�O�~k������Q�`�#�CP���e"��d0E��;�CH��޸w��H	��IgĈ
:s*q:ץ˳ST�R�$��$/��>zs���BFem�G`����fL��gX�� �%��BAjk� �_>��ˊ)�HfL�2͛i�Hq��sE���x��_���]
#��RV�)��ʅ�3tC��2�)j�����azu�n�(�iV�	GA���4�*H�e�j!�P�ΙZ�yh$P�/wh/��0�HQ��cH�\D4��ONvCL���!�Lӻ�,\���R�PE��Vh�Ԝ�ȺC5�G���3)tЍ�jux���Ve|a�8�"�bSLo1�K+ӽ,Ĭd��1�Z��R+.2ڞ�!S0�U�A[H�FM�������G!�C
��X~4$��#B�QL���S���2�r��ҧ���e|�����b�lSJ����n�/)֯e�vE�9ʑL-i�"�燏��m���sm���H�	��z�Y){}�z�ҳ�fK<���+��1b^f%V~�Tlh�U,0�@,�Fu�����ae��A}0�aq�W�lfF f��U1[a�wLh�#D���nC�k���}��9�@���{������9��WΜ/!��M<* $n�G���K	JC�)�>�ɹ���x�TT��Y��%��Q	+c^��C}�x��(��`<� frմMY��<���Q�)�9?��B=ME�[�/�;D��/����l�CKQao���֮�I!�X�q3��h�`��]=��㌳U9��v��~4���	d�0BQL��t�eH)���$u��ʕ�C���LՉ9�q}�5e�{���d[,U�ϸ�J��Ƽ����@�2�:�[T"��S� L73�tE=,U��vbE� ��T�3K��%	�k�ݕ�n H��661��}qtL9���4��Ƃ���I��@�@H�jZ���}Y���E!�.CAŰ����;c/$j(��š�5>��$E eL� �G=R1
��*���e�7u�$B�G�{��6#���$g�P��-�CD*�`��Պk}'[�OA[5�s��W��\��H�J$�;�����&�/*֙.��`��H�^�M�_о��9��KZZ�M`��%s�h)P�y��!�MuÜ�Y#Y� �9�%C�<������9��p0`$W3iF��#S!M�4����Z0�0�S&�:1$༂D���
[�j�i�a]�p���崫�!u���xQFch����fŹ^�is�2�d����K�.�p�!2bH@