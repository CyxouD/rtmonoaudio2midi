BZh91AY&SY�Ÿ �_�px����߰����`_�� lp@��A$��6Ry��jx��6��x�i�2`A�~�� � @   h�$�A�d 4i�A� 4`�1 �&	�!��L��`�1 �&	�!��L����4�<��Ҟ�F� i� �BFG�΄�f$M ��X O����HG���*��0l��0��d��`�b0EX�8���Vk��vz�c�HF����Ǳ����,�bi�Nh�hq��B<�A���-dr�2C6W,X���c��Gy&a�Δ�����@�V� `/� �i�T�B��������=t���ҶR�w;+( �����,��	�r�L�Q&T��aH�J,�)D�R�
Yv��6�J-���^���tw%ߊb��PŶ6F$;��4+YT����ڈ���Zh�M��2ы����B�al3���&�5z�m)L����Gaf�Jl��31h�t��������d["0FQeI�Gv��KS&�i���TKm!�a��d :�g�zJjv�L��ǲL�H�0TcYz�P�IwhS�C�8�|�E͎�E�l��-tж�S)Y�æ �4�CT�-����t��E1/C#%��w"/M8blKp�s눯K��~�|C��	�9$� LD�� Qz�R+:+��!H�M(!U��e^A1��Ԕ�D�Cb�?VC�8�	ix0��3��!d���OmnhBld̙�����/lq���V��������@�û���[��|eF�f��3͕J$#}7yn�Յ$!��a�3@�|d\��t�<h��O�Z~5�R�Z�b�J6�����R��a!f��O@��CeЬ�J^��B�'�4ȏ�IO&;���,�)zĄI�.[@�)j*�i$Sx��o٢f)������=>�+�Gfv�����M��[�R�P�^��g�p1-��I�\`��:dҐ4�K��pO�
�LW$v�ւ� D��9fW~��X��/����^�D�z�Jオ��w�����@���ϱ0i!���$�)�ګ��xP~��u$�d\�;2������1K{��B��1�B"˕��z����~"Xx���g>KLք�$#ǹw�����w>w(D��,CAɬ��EBZƘ�i��u%�Hj^�i$"`2�ԓ�g��D�u5gV�("a��L�v^%D��T��`Off�r	�$#6�D���P�/�=9��bj�c�c�OAC5ns[Xl�f�������)�"��ǩ�L��u��~a!��YT�|Ko�ͻ���IdS���PGL��"`�g�a�z�~�e���م��ȕ�\՗D��1*p�C����!�[����Y
V �9�Zt�|^�1{Ƚ����&�\ǿZ_�_�@�W\��S���"����d�����dn1(�b_�v����$Zɒ3P�l!?�]��BB�c�