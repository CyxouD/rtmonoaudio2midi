BZh91AY&SY��NU �߀Px����߰����`o�Mƀ�D�(*D�AS�=�g�h��ODdzA��=L�P�~M*� �� 2i�&M  �4���4��!�d2�2b`b0#L1&L0挘� ���F	� �"&�4M�S�OQ=���L� ڙ4�;t$�&a"D�:@�)%3�x�� o��,��  �0�����I��1�w0��V���]>�X� �V����@u:n"�W�_#��Y�9(;���Q���b�P���  �v �! ����4�/%�,(��j2�ln�J��6]��8�8Xa�z��D�2�Z\w ��9HP������7ͯ���� 3�w�:4u��NW��Z,���_�u�{�KvB"$�ҟ�1p�L[�����jRSEӸ}k�h �l��3���dRq�%;�-{b)ӶB�Hj�~�ݭqL��CD5�(e}ε�HR�w4�uk�R�X����8fhҹ���qI�9sa��옾9Cr]�k�6EE�X���NY��+�++@�`�U�r*6����mc���� \;;MJ�}��c�S�ܸ�a��{Qf-k����PKE� �)���r��?G&�;Ta�܊`�j��ǧ��q҃���o!�� �i�6Vr\�MF���E�qU*l��3�K��]���W�׃�,cB��o�	�L��V�Z���.�,�XQ���ʶ�Lɢ��wvDuLX�8����ź�����Zʚ���7��D���l���X��N��A4mc&�|sEk�]`�{Ò�s���E�#q�d�9Ż��l�?o��{f����m��4 A7zzT�%/o���Ԭ��.d��E�k�Y hL`��K��E�>R�,� E"�!E"@ b����K���X0�a{U�|�HfB
���k6��3���~}�t���s����wl�?��nj�b+��dS��E*  w`����V)P 3IӅ�7���RG\��t���ǟ�y��� 9��;þͯ�>Į�^� �Bg^}Bj�V�O2�&J_�x��9�dy�$�x����gGJ�ۇ� ��g�vc����:e"���� ȃ��]��f�(ȟ���(U�)��ڝ�dҭB�i���@�#BR�,J�AGX:V�2���u���F�Ґ �]Ϛfx�f��i.�����RMM
e �� �[9�㛝��M��� B	��hU��)�f	�i&���� ��m09������f���P�U���3� Z���0�A���A��<(�Zc���X\(2A�Hn �ڽ g�}v<��s�b> ��rk(��N��4ZH̢w�B@@��U}�k$E e�T� �|#}R2��*��B\�!ܢY��E� U��`Oon�b9@ � �%�y�r��)�UCק�5�%�o�AL�;�{/�fe��-ga۽+K ɏP#�2_����5�� .�q�,{����}�U�r%�q�j
������B(�<7�����[��{�
�"o��
ˮ���K�i|�  �f����g)�l�Ki�y�~��_A�HX�&�l��V��IrX�)gAv�UFmf��� iG��U�/��m��,BF֚EՏ����.�p�!c�