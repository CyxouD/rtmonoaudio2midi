BZh91AY&SYM�j� p߀Px����߰����`ώ&��� /��%@�DѠ�h��hh$��Q�<��6�4M�5=4��M �i�  ��OP�       T�QL�T 4  b4  �101��&$D)�S)�Oj��e 4����Q�p	�$H �I9��h���eF]�`��5>R�@�D�A�`�1�oa"�0k�Z���͒L�ŉg��Nc��+��-L�6+T��*=z�����6!���B�")�.&��)�E�$#UU!	�:(K3Oܘ>p�%�f�Hʚt�ǫ��0H�s�%r3µ�oA�*���jꔒH�/,��������?�ʋ��mح�[�lE�P.����Kɳ�Б��I�҈h�](`�%�����2�Bq�T0o�q�Z�B�g�z�Љ�Px4i�Ȋ���$e�v��Pj�	�|�͂�v���>��$]��Z,=�k��ͪX�(��Tj�ډ��*A��̤P��jk]KE���2�l�O��Apy���AY�C�8@QI�a�E�A㈡X׀澖�h;�pD=	��>�#1Th��u���U��D[��h�L�mg7L<Ak݇�f��D�"(GN�g�x�*E4Xl׷��4!�떭3�`�$DL�-FR�����{����,=e�M�:�j��F�U�Dmk�ˉ{�Tp�����vy\��6�2��R����9
�Iw6*A����V!���ESW\gp�,���7-*ⅺ�5�Y�e2wzN��˲7j%��Yې]��号�G\���!X�Զ~��:mv���CƳ
���]��z�'J�Z�8�<�:ұ6�M]J�d��d�Wsx�-�h`��tajw��c �=x1,� :@ I�A�o:�4J_w����,�+�1vK;�0�Av�B11d �c1��(�������F���1oasD��9N�2`�(o-r@� ,�b�����7a��דy��c���]��S����t�~�=�4��U�ǝSl�:�*�����Wb@��(�y	yJCn����h�a������e Ʊv诀p�}������ n������z���U)�S�?��a�m�?����.Կ�p 8��@ ��.,f�i�*3�"��m5P��tE|v8�?!,(��E�3�ч�˷V�i-B��Mu�� .Y�X�!D��N��L􂛠�:�Ga�۠���% ��rܚ�4�_�i^H2�f��M�3͊��� ��^���GL�Ў�/յ0b*�"���m��A�q���%.<� ���v��k��2|a���丯�]u�s�cc�����Qϟ~�Q�h�����]FV z�WR�d#��dw��a��T\��a(�	���i#ID�NI �5?}�$E eL� �����EwSy��$ �(�lw^%�U��'�۠�F��}D�6��V)5IN���8�ؚx�z
K��gV��:V6H��&�m���#�@�iԸ4ЙG��`��!W��c�п6Y�����q%�;�Yj1��״�B(�>'5,�o�7F��E4o��NR:�J�EA��L<��ѓ�tZ�eGUs*�K!M�2	Uu��̓�֎�G��85$KP��5RӰ��%��C9���&�EN�[a�3�����Z�3��sَ�9"�L���۳�
��H�
	�mQ@