BZh91AY&SY���q _�px����߰����P裀�Ė��.�	$�Q��O ��FM4��P4��� ID�Ѵ�h b`��%2"ji  Ѧ�hh�4  �=@8ɓ&# &L �# C �"d��SУ�#)��&�jh  @Lߝ$,$A$�9 EI$ߓ�� ����) H � 
�����I�Q����4�0��^�v7` ��~�(�}&B�����%{�)�bc[8����,�RJe���?΍t�����$Fw�О��F�H���i+���\Ǘ�x%d�  ���:}ے���a����V�����Zv�,�`ހ؁��_���e"U%S#T�1�SUSո�r��85�Qrv)Շ^��Tfʝ�x��<N�O"��j4�m��fC�).X�E�A�EU{�Wt`�&EJҰJ�����g!h�l[��Q���3˔-1��@k:3�BS�V����XsĄ�Ut�f�=@0�X�Ö0e�J��iD�C"��+$A�:1*TR.`�.�pqN���a��f��1��˼3BI;Pi�dE�d4,g_@ja���A%�V���;V%YcNy��|~��m������I$�( ɿ��&#��U�*��n�q7kA�$��#B�F�1(.��"$׹� �"� iw�Q_C���aQ�L��Z�VC0�Sbl`kw��*w�����fíz)��b�	f���w�������vPXy��א��YԀ~�����ƀ+�,��#ͫ��#ƌɽk��x�mN�!���fׇPuU���B����hl ?����'y����}�M+z�%2y�a��?��M��Ҽ.΀�^u�����|#@���F��G0������=��/�9۷	J	ܘ)���/�A�5q+�R��C�<�p4.�2L�$*�$Ι\,�p�郈��`XY$ W���3�zV~��]�M�$�%�.Ȩ��  �Yжp�\�?�4l� zpl�P�5Qr������#�=+��&��!.�MZ����*o�6@ ��fk^�O�@n��}^�H�.�8͚��\/d�`յt�����m}�(D����!��HU��,F��I�4�Jք�Ի+�!��' �xF�2
�4�b�IA%EfgU�( ��A=��Q� . <�(9�c,5Bz�=>2�t������������6�kH���t�ؕd� M�hE{�	�'bH B������W�f^(֭Ja�%@�1�;F9��;DÄ́�w��j�@i�u��q��2�t�c]�U!
�`� � �z�z�r��*�`9�+,��n���t�<)I���E�Լ��Y3<�]�k�QLU����@vM ��Q�YV[�ͦM��	ZiW�ݬ��_�w$S�	*�w