BZh91AY&SYz8]� ߀px����߰����PM�;Dn(����	$# �H�z'��4'��44�cA��2d��CM     BBMOE�4i�M @ z����a2dɑ��4�# C �$Ě�S�COQ�2Mz&�������� ��Ԑa"	 ��E	 �x��N�����f6�	5}���_�F��ch�a"�-k��gۍ�^	-4�&~~�A�ｼ��w['w+-!ŇD�\Q�И���G��G6�n�Jѫ3<k����8P�͆�|%��q{:b���I$L� �]YU:=��]��M�G��ٽG�ȼN̛�U�ς� ���٬'���L�D�0�5����4F�qhsQRTզ�#�V��o:����a�Eڂ��U�5t����fD�"�JX��n7$���^�鱢B�[���*�US�)
�c,t�i5��U�SX�n��2�.?f�7��m���F�m�BP�c��U�)/O'n�+^���)�2_6�5L&uLi1�f��P#d��M.fW��d��*0����!3%UN+k�]�z�F�x���p����Ǘ�������i�w�m�E�}�^���=��.ۿ�����!&)���D	��&�d�ͮ����-��ǥ�t3Ж��ӿ�5}��!s�����%��]�D�87�o�ar&J������Q�(��7n�ں4�@s����-��j�h2t�)�($O�'��]��!��D��s����W��*�g=ģ�ϙ���q۠�]�Ҏ1d1VTo�J��{�u�Y�
���5�Sj@���<8�]A�˩�OOzf�����QS/ �$��[5'�o�gي`d$�����	#l�����A2OKED�pͨ��c����1ch��>�tq�kM %5Y�fk����&�={��]eRek�HF�K׽q�#��ol��D��4T��B�f�Y��+"0,N��h�r尡�5*N9b;7H�Z��N]VUe	A
΋�yJ+��ؽR��,A-|�Pz2�Z(e
�LΟ��n�gOAQ{�ܗ�d32��GY��lJ�c�[���$�Z��yA(S夨m�GMt�e
�fūj��N�>�� q��,��-~/������5�RXV4 $P�~������q��4o��A��'V�T���:RI���D������a��@�׺�r��'�EI��㗕����ኝYooY6j�H��H�y^ ��.�p� �p�(