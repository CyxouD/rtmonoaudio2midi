BZh91AY&SY��� �_�Px����߰����P�8� 㸪�F&���	�M5E0ʙ��M0�mjz J�       ����I����6�� 4�b@i��2b`b0#L1&L0D�LT�
2��S@4�4�4�+�V�V�)`"�����w�|������.� %ʌi�:�e(n�0 %��: R)l�Ͼ�z��eTuJ|v%�� 1t����x��ZU �E@hi�i��66�6��_�ĝwm���P��3�c����̙�&Lag�d�DV�vUq��j�g���{���4h�|�e=��bm��9�m˧��|�9Ѓ�.�c��ONt�RJMP���-�-�:[�eF�� N�"i����;T�����1٨��FK�8^�KFI��b�6R
%z��c6:��I(�&�AyYaV�S���h�GXF�AU�[1ʙALU�ag2�.�څLVWU�f�"G���� Ӏ]�tuM��	��u���w��xA*�	j��.�M"��#��1�m&���4����:�����ڽgllm�[m���p�
�bR�r몵+;b0d��"�[�WhF��D�������U��a$�ed��쁈�Cd�]��.`_]�9` �ح��s�'.�r��.:n�z�)Zޟ�p����,����g����E��Zvȳ�N
i!{���}~�W^LUP�i�G<s��#�:5��tU�q�s-f6 �OE�p��>��Q��$���IG����t�Z���<~�+���G�v�D��k�1�h9>�F��CNBXe�-N��0��cɂ���k�s��������U��[�#D��>,���K�t���1(h���bM%2F�$u���H)��26�<+%$'9�;�S7�[�r�ц(�٭�L�
�*�P��|�!RF�A����
u�w ��@�*�/NKs6���$;�Kɂ�4���0O���1kÆ��b�,o��`�g��{�3��#�O>��>�7V�pRka :B��u�^`/r1n�M��"����,CA�J-���7Ƙ�i#ID�M�  MOE��@U����qb���m4PD���g��0 I� ����{,/F���$��H9o�\(o�|"���:Ü��`����9��ٸfŃ$j(�&�ǩn�"�3��	��g����7�hT'*9P�W���j<��J��٭����: �i��#<��^S��AJy�T���lT.�D�C�쵱�HT�HTYl)�Ԣ��r|���u�ΐ��b�6�Ә�(�m����i�Q^�u3�n�"�T�܌th�|lrH�#��t/ۿ���E3�)Ð��¯�]��BC��� 