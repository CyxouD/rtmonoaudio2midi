BZh91AY&SY���U D߀Px����߰����`_5��$��i�h4Q�S�'��1F�z��i����!�@���0       sFLL LFi�#ɀFѓ �`A��2`�4d���`F�b0L�`�B)�d��I�<��(��4 `�J���H,Ċ$�(HH� G�D��{W���eF]�`����a��D�Ou�d0E��<CH���<u���p�,�`���ѽו�e�����6��<���tX�O`�LȇrC֑QJ�+O��OA���e)*J妽lq�p��	�35��hЧ;����R�2$%�\$�{�g.x�00]��+m�:O'Q��gb��˪��#�k��n�o��j8�#��5T2�kiMT�g+������Pور;h3�Sv�5�0����^?��~n8o�HFϭб�K�T����fL� i��6�2��0��cq��M��=�EiH���3P�,��}���fƃ��8]�i�J�u��r��L�*t���n��8l ��uP[U)J� �Sz+5��&ԌG(�2S*0��K3A�|7*ݢ�pB��i[f�m����m7�u�^�)k����S��ơ��!@FǤ.+�����^F� �߱��`� �	�6�>D����W�gTE�,��ׂ�?�	hR4�0�`����&���VA�H8�4�P]�*i���}P��a�U�͌�bI6���K���_��-�qW��-s����6���>>���iNVS�,4�U���  �Ww���*��@Ĥ>�/q�M����c�^����z�f��U}.p�2���}����N� �93��X��[w�ز�ER�آI��w�)l�[���ͽ(#�_�-�[P�/�u�fzD�D����f{��_Ll�p�%'h�y��Q���|<1�d�7�}�bc� `��B�Jd떔�N��M�mxIpvЎ&G�QQ���t�ݱ3^%��5�#P�l�9�Sz̋e����w���<�B#t�����L+�C@ګ�-nUn]��XClA�YI]8�(2c�bы�9�Н+]��W3h
��cc�}����N>�3J;X��[#$�fV��
܋瑩���P2 uE�h3�QUT�����3(��š�5?��$E eL� �8GER1
��*��EHA6Q,�w^�����pOof�b=  ����;�z
��O4����!������Rͅ�o^��б��I�;�ذ��`���p.8���{�A
�כ�_��d}\�U�lK@v�k1����)P��?~���7W��pņ��fy�_&�xc�ᄬzqx���X-��|��h͐���B�<�a�z9���#	�ĢE��~�>kJ��9)�ud�����`��m�o���Ch��Un�?�Nyl�$Zɒ.�v�!/���)�t�¨