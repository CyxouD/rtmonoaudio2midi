BZh91AY&SY�߀G #߀Px����߰����P��7�q�ږ3IBIhA4�OML�e=G�h��&�hbO@	R    h   	������ѡ���M2h 44d���`F�b0L�`�E3)�)�F��=&��4Ѡ�4@*z�H�$A @�RI��N�;������Y��.	C�?4��BT"�6� �*a6�l^.�*Z	���Ȗ~���u�"�^S�μJقo1N����u�"ũ��AbO��{Lnv���3r����J@���w���K����ua	��@�_��i�C`×��M:z���5�ŉ4kAK�u�8��a�3?�����u�6���-�a�$ N�"h0?�F�=o�\!w���P��u�kH��[7�dTٶJ^�C�v���j�wFV"QFK�Xu&�
��Q�E����͒�����%	�'[�St�K%��)Ĩ���� �\T�n��l���OH�J�r\g���Q�4���t�*ZV�be�V�Xg������Q$66��m�	A7�w��7?�*Ӫ"�k��ˬ5	��͆d����@�w�h��)�"a�,�	\�,f����xV0�a6��X<�m	;k���ˬ��N���p[�>��	]��W���|�����i��U�M�9�+�FU H��}����ء!�ie&혎�\^���T����núE�Ƅ$eY9,�'n����A�!�$u��_�P�cS�[�Z�Ћ�neN�-գq�H���X�݂��b��G�%֗�qCQ�pJE��+ǟ��SJaod�7\G/(�T��613��e�gՃF'MU��;�+m�5�D�X�D��N���Up�pv�G�i���"	6�ze��t�:�2�o��)�ҒjhS(/��A{�#���4�_Ę	��l��hQ�9��W�A�|��m���a0[ri(3�&2tF,n Ò�X�ϒ6�`$F�Xflok�,���9�p�e���V����k�ɤ%�	::�ނ2w\t=N0F`�{�!��J1J��4Ƌ����94	@���g$E �)N�0��6���S��\�!�D�K���
�<��z�1� $g�6���ː�(r­q>r�:$a���*1�ͣ=�0s,���r:M��IN�$<���2/�m��D�tK4���+�T{8�cJȕA�JЋ@�6"�3Xuj4���	0U�U�H)�Dʂ�эje�J-�A"%f�nx�3�H�ۊ��Ɗ�^�(ȁp���y�s��!9�	 �fH�����a�@�k��r츚�:�����pBEl��������Ͱ�FM4�[Ho�)�rE8P��߀G