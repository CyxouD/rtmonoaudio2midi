BZh91AY&SY�(�� �_�Px����߰����`�-���R��$�L�	���S�=S�ޔz��=����ԡF���#� L�0&&�	�&L�&	���MSM4�ѵ=M �  �	���dɓ#	�i�F& �$=2j�zj~�6�&'��d�@��o�䢛{��SX)�
A�B�i�}����n!�	?�D�@��1T>��g	�E3��|��ݿf� ���^��=�`J�J���TF�Y�T��؀�i�(	8����,&�ZN&)n��ˬ|[A(�u�K�O�3n�Bs���9��y�v��1.�P�����m���|�M0��d��}>Vtts=7�����pi��s��B�rr�F�{�o͊-Li�U�i�L�~v�#y�A�����U͗C~� 'bD��n@l(�a�����@LȗK��5��KhM�K�:mG�x�:i��2^/&���j��榡{���2��#��-���QO��5h��{5w�&N��H"2�`�R�,��Zi02"�]�t�m��[�Q����w:���@��B̲��/���I��Ռ�m�T/MX�P�1ݴ�I:z,�K5,S���`w=�fN���c4u�AܙJ�.-4N��
,�c����s�!6Q6�1Gf;�΋�|�����j����������$Z	$�A1��c�y��QȚ������-3tՐ!^�^$1D�*(Q�(b?�F�6V�V���7m�Mԫ`��6Q�C�)G�'|g.�r�ν8���]R���c	���O/G����x��/9S����b�t���k���e���1d��W�
����wDxѡG���w�Ď��ƴ������97���h��� ���&v��W%81لTMX�"D�f���ƴy��y�z���ƫ�Y�ĄK�/6Z4Ѭ��2�6�~�ױIq�j�����]p�f�$���Aw�19?;�Nj��?H8mL	̀Ԁb�er�3x,���0�lO!Y��Dax��>�ZoL_Y.E���1*v��Lً
��T����B+#�2�.��@s�Ӗ����R߁�SǟK�O �<�#�[����?AC9V�ǙQ�1{h�0r�X�ƠHDi��a�����vDs��p���c-��3[��Gf�"X�}<3�E'T��<�L1;d��,tÂ��&vW9�f^�@hc~�7& �F�����rS�:�f�Y:U��]��W~h�b�R�;l�6�6�#!D�z�Aտ�C|)�!��}�@�3w{��`��9���!�=�l���Y�y�k��
$᳊'c�<����쫌�#��'��4퍋�٨fa�$��g����9�>!�k�M�ݓ��`�=�*��gj���Sl�&<�ʻ��!a!��4��b�/a��\4
���u�k���Ǆ�pn �U�j�/Ejۼ����r��Ur����y��A߅D�"zΗ-!����r�����k���)���"�(Hi�[΀