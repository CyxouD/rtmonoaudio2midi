BZh91AY&SY�lk �߀Px����߰����`	�|�N�a   �8��Dl2BI��	��L
<S�hi���2S؀�J `M F�F� �101��&5?DR�h4�4ɣ d��M "�F�����   ��h$D$j��?BDڠ�H�����=AzqUr��  �'U$
p$��	��AWO:Y� �a�g�G�H �`�1�{CH�5�Ҹ}=9�@�\e;o%��t�u��e�F���L���	��	2� �GWW*;t趖0�$�!G	r`M
�v����%Ɉ;�*�bJUn�U�*)EX��j��L6�����i��6�BFl�D1Ǜ��PHǨ��eU�����9�S�R@�1xfm��yv�2�fO9e��pڳQ��LE��^wle���_me���a�cʛ��++��A;w�N<�5'`�H�1����1\:h�WY�x�r�Tؖ #F�sC?��u���� �.�ۤպ̑��D��1�1YHs���wV+*�F�k%c^Qw������6&�yY�,`�W��Ǒi�5f(g&����e.BX�w�F�kIE�fY4�]ݝ�Ɩ�5����fD�6�l��6p��!�8�:�7G,����2�EQC.
�G@�=\�B�EI��2n��Q�S�ۙ^�TLwPzg��9�K:ś�� �8�Vj99�)Ŵ�S��]�߶/Э9:�s#˭�VE�g="�N��F�n$�݊�2 �vrj����F��'!)���U���>-�oL��flm��)�Ԣ�HE���X4�U
��U�R޽R�9Vi�f[�f�:�7o!ȹ���lЈ��V��X�e� сV]ص���躛�p�c*�%���;����9e
gwo��-(u����Bo�k�/$�ı:\t���s����t�Au(��nރ�t.}�+*����
�ĲI3A]��=L���(�U���'�)�z�<�L�Ȏ�Cpe��uT32!V!�ˑ�R����Z0�۞�����u
H�ؚ$�ۤ�%�˘x�K�}3�c�ȚuX:WEb�=9�&���C:�+���j� ����ȍdE8ݰ9�@!��E���jSh!��e�Dz�ړ�3*�͡���,+����!v2���R�ug+ͅp��x�n$U�4ƾ�)�Ρm��tBvK�H$s�D����¸�~f;�vcA�>_#\)t*��?"���.E�( 	�je�������v�^���;�vQ��7�	y�a��^P��!%&����ZCh؃Y��I&.l.k7G}��at�W�6�����3Fj��Ƿ��_<���f��p�vxJ�#��	W���������+Ņ?Y_y��V�.Q@�]�h��~�YjBI1)���'&ߧT��:jJ^�˴ߴ�D���!$�X=�,���xz�\Ƞ-��AW	$"$���nǾ���P�:�LM�N�{�߭1���VZ� ��@�+�AV��c=C@���G#�&�'��%�{�����q�%�(��{��Ǿl�~�zn�KP��ߝ}�}�$��	iKB2@(�;��iҹI� �,���drԨҫR�$��[��3�"��1<��9��"yP�P^\�J�kxB=S�B=8���S*�R���ձ��X���I[�g(1�4(L`�'3�V؃W$֭���̂����35�m�7,ßGF٥V4i�1}��Q��@P$�FE�|�n�u�f��|\�(�QrĢ�T'p�-$tN�� &���DPT���T���EwSy��$ ��SA�<� ��h	[�P1f���g ��Ij�^A�^�C\)�0ztzF�鉫��OAIk��mݠfb��0�Gi�M�(��@�M��`�����ŷ``́$���;�;?�����ɪi+R�7EW|'a��p�7c!0: �a��f���iٍO+�D�F�V��.�*���X�Ǿ�K&�$���T��UGC!M�6��)�n:$�F#��d'�l���Z��.���&r�g/X��r2Zg�����?�V��뻲[;�;i�H�3��ܑN$a��