BZh91AY&SY0Q u_�Px����߰����`Ϟu�� �Q UIɡ��i��6��h򁚍22S�@)I�b�� �	�=@ѓ �`A��2`�L�*d����4   �101��&$DhO)���z�)�H���h �&��tN�jBH�!$I	R�B�x�y�����;*2�T&���/��	b0E��90��f5��Z}9c��v�������0��3�^�N��R�(E'$�:t���B$E�)�t�$�`�F�.�v.���_���u����-@���z�
�S]���&�xe��,�S{��l;9I"�H��}x��ܾ�ϻ�f?/쭷���Z��͸�,����}#�P�"�40o�6t�&�ō��W.��!Pme��I��2��i�����r�K�`�ˁ��&�,@v��z�5W@M-���d�,�	�(Be�Z��f�'ahv��&���vP�P ��C��(����۷B>�}�iS�3��A>#�`A��1G]�\��8�fS�&��;MS����(����Iub�+F�g��RmO(u��6�!A�bv��T�X�ϲd��p�6���3��b�p��tZW�BV�|��DNTrL2�f��^���0v�\��oN�*݅L�hx�LEʜ��85�ʃ3D�����X"خ�^ls�4�]���;����Aծw	61�ݮiFx���燳'>1|�	��I �`x���fǇv�!�Ғ�IDI�ȁR}%�cP�b$iaŤg�ġ��жD\&.L.l�����Z�]0���,��$3$�j���ow\a��%.�xor�w���߮"�^ώOώ�r�x��+�5@�E2Q}���p%{&Re3o��_��Ǎ=EOP�[Oq���xe�s���y��_�|I^(�4hl/1���6	�9��6���'J����˜�B=ME�s���L���@��.[X�2u����k���$=�W9�6	Fd�5�}*��,�s+P�n4͞�@�X)h���i$v� ӥp�AM �i֏I�ߴ��VA��[�$̵�/b�l}�"Sy��R����p@���4�DRDZ����
e@w�
�#KpV���yOR߬����j8n?���3k�uН�+�g^c�
��1��9~��*�:�����٭s@j8L$	3�/.+�hF��s��s�b>�uE�h9�(�*�NcLh���Q;���x�eW۫2DP\�Jp�B4�F�`���o4PD�e���XB
����}^����g� ���%�M�5Z'^�X��9v;�=��&}݃a�4��#�;������@#Ja���i� ւ�G=���C-�:����ZÎ �@ �7hR���oa�L��x�Ulk>�(G<⤨|h���k�(3�cc� Z� V�4!�Gn+*&2Up �+��!�%2l��� 	�(�l�@�U�I�)�/���3�qE�
.F;��87L�
���jx19^�s9�Y2Fj�t�	�ܑN$��@