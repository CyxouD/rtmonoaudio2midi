BZh91AY&SY@��� �_�Px����������P�9n ��zsX��$�F�����RzO%=&�i�44 �d��1I@&� 	�р DA�<��z�P4  @"���i=FL���ɂ2d�@�4�I�z&�#��6S�I�� hh@*�����)b�4U*�AgQ���^�����]@O�+@��2uX"��H�`R)t1ա˻��`����ϼtپW��f�$�K���-�R����t�8�p��	��9I��%9߇j�l�UU��Uc�r۷�~4a`*�32m�~+ׯ���]���M���z����7>�ls�DGA�K�b�p������jZ&��y`�i�~T���\kC	 ��"�H�v�Ml�|��r��˖�g*4u%����A3�1b�rp5����H:��&���:�_W����[k@xh����C��U �>i2BhB�Ƣ�u���40��U�K	�	�2�R@�)������b�4=۫�	�a�m���p$.ѻ��ޥ��#[y6ҡ	�f�E}<�o��m���3m���%n���bR��⪽+<Qd�����l|�%�3���g��UV��#)�H�$�]�Z`���,X\a�Uܵ�� M�hf����G���y�4�v3l�Q�q���r�Q��4�׊��j@��'����߂[�Y"����A]�Ψ�6Y��������b����+�C���x��,!�$��]$J<�Q��r�MoD��<�Wr��F�Ѧ���^1��@w-�z�%/j_V5�4�:�p�"8�듮����r�����wWP�Qɦ���4��3��0��f�j�r�[6�
�
�I.��#�	�k��)6A`�/Ncx�c0����"��d�.�dr������JoQ�l�VT_���Į����؟��'��02Ozpms=jO�3�j��q��z�ҝ��yg����BGQ�b�xr��V�:��� 	(١�a������ϫ�����Ӌe�
#�C�������s^w�,����A�!��$W��:�c-$fQ;�@���o�"(*`�8z�H�X*'x��ĔrL�e��u�,!%
�;�������$��)A˳|�P�<1�?t��=.Э�L��Ï!�<JL��r:�#�4�X@Vg�B'y�eN��	����wYq׸���8ְJ�㒆�3A'�E�"� ����F��0[��=�T�8����T��V5��UsP	)0$�e�.i֢��r}#���B��%Pa:�mC�!�JN�(�mX%ޭY� h�譜�+�(�R��Ox�l���t�C�.z�i�����&�6l�c����"�(H YE߀