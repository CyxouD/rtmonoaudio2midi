BZh91AY&SYן� ߀Px����߰����`���z .\����i?!��ੵ==Q�=��L�4��Pj�d%&���0���209�&& &#4���d�#jDj'�4 � ��  9�&& &#4���d�#��=�Ȧzd�<SmQ�#F���mC$RI�� )0�$�t$,H@�`%G��/1	���Yv�,!!�a�K��@�"�m�CH��޸}�����WD���.���ǌ�����j�"��J3��2y���Ә-.�g��w�KC�JtJhG��c��`�z��p���͎>NYA#4fz�es4�Pa��­�BH+\��}؆�r�]�&!!�a����}���r���ͩ��j��4`�^�Дp6F�r�0�(D���^�߄�pI3�D.�z`-��n���(���I��8�5!��آ>Ҹ1��-��U�C ,�\!1Dtn64j�T	�̌ZZ�Y:�CF(ش�Xe�.e�"����4�\�9���>�蹎��%�%n@�Rq��,!��;u�Cx��Q<,�[a��J/���\E=ӆ�M���ql*^�+�C�ʃe��wl],;�0Fu�l�����2d�%�>RD�ԋѫniK�WOMO�q�]N��DLI�m{�c Hc���<��.��5�A��s�
�Q�u�uS�N��7�By�0��j��'e�L�ږD���+b�d�f�rF�rs���g.�x 	��(R��-e&��ߩ^��؋2Y�Z��"�<T��Ra�"�Ҡ�����)hKLE�$1rab�\D�dðJ�J����"`�mXX+Kأ�r�'*��ӛ��r����	]堯���Bx��O���H�ʬ�7ȳn*��$t�W��̫T��*����S񤣆������+��Σ����b)	�[���3/�z�^�L62�$}�@��Ә��s}uoZ2"��w����)G���f��u�@w��.�y�u�D��ҋ��F�Ap��$A։���Ϙ���R�1+'��|���P�����V>q�-�`��"��N��L�:�:�$p18�,1�	:s�ԙ�#�J�A��[G�dJoY�l�VT��BF%y�w�����b`�&TC�Su�j�ޠ������ �Ud�r�y�Ӝh����-n��THX�_n��t�+��cc�{�>�|�D��ƹaɛ�,�16L Bg�BG�r�8GC���9�P2�uE�h9��FU'X�/$fQ;�I�x���Y"(/��Q8~P��$XX*+����!�D�c��,$$:��@���ѠBE�6q$����b��m��~'Xs�����V͕ݽ�{5���gd����N޴�,bV\S%��\{X5�SƘRxt�'v:�޽�V�%`q��0�@q�с�֞����D�w�äT���h'[J�짧 ��c~<�m�$b�$[��'����U.A�:Y�C^�r}$a�!p;�S`�y@�V-����x�΃]�ڤ��Ӑ���R,��iTI�8���A���s&H�h���_�.�p� !�?�