BZh91AY&SYb(�� =߀Px����߰����`_.w      =ÊB��	�S�)�$�T�S#j4Ѡ�F����J� �     �iT�#C&&	��hi�M4�0!���b�F@��  4挘� ���F	� �$@�5���ɦM56�&OSA� ��4����w( 0R�*�@�9� ��-|�����|�86�0$�AT�@�<���;	�$N���r�Yp��$	$f���{�	�8�4t������d� ���A��XGSu��	.	Y��ڛ�V�*�+,�E*q��,lM���ZUGQ�RIBaB�� U6�*b"#M�-M0L�3(�`&�!��ɂ8��`��਼gͪ�$�[Bj	e,��H�Po�,8@�\(�
�vE-,G~�_�K�3��T&�/W���%:iE�la�[SJv��C�0���㎶T�=����y�b
����������ȰhS�y&�`�la�c�0 �3�(���n���%��=.��陵o������`L���{�r�|u�Sj�
c&[)�aF���J!UR�7��ډ����$�bX栅;v�w1�D�╷S��vj�b���b.����w"�'[yǿ��]�O�����5�Ǥd�h��_�G��G
����>i+��C��	���Ӥ1/R��"=���a��$D�a/F�B#O��+�a��9�'��1y�"9x��$F�$�>Aj�qQJl��$���(@YA�����H�2�����di�	�A�Am'd\Fv�ZM<��^D��`���E������	��"k��8� ��y�j(Ud�H˦&��^�Z����	�Ɇt�E�u�	hY$Ok�F�6�8��)5���F*/f8d]`�XV�:�W#4�d^n:f1���v�qLEe&�F��Nqp0.�,�uzE�^o��;�ރ��Uk��U���<�. �ZM����4���Wg,�����C�v�*���.�z(NGC�`�)�"ž��Ą�2E`I�>�s��eQdF�7���Gf��Q��^'1V��LA��DlyU�4;�QX#�1�m9��&0��m�
�"�˛��J�	-n!l�p��,��TG)�v�3�ᣪ�s��rB�u��U��MF+�{Y���43����2�Y�<Wi��w�;���Y6�v"�t�^tk/C��}�d#hَ�.��b�N<B�/n����P����	��7�G&* ٍ�w�&��eś�VHA�v�b�7�=3���2�WF��1/L�(�έ
N[s�'�̽��t��iJ����R[���NNaWt�c��<�հ�o�VIq
&��GB��I"�V��G*Z����'��&���l����M�*�Xc�=��Hځ7D�<عd.��c�����a\�Qӓc6P���Z���ūBt]�Wʱz=��߮"M��jj��vr�3Y�; ��^3��j�PrO�V9v�S�kj�	�q1�2�ϵ8:l�Ò4`Q��s�]r�wy#��ʨy\2g3] �s����M����y9�x�9�io�Q
�nBQ�;QW%�G�x���n�s�L��"Zy��������n0eX'�Uf�]Q�"���SH!D�$XE^Z9}Qb��yLb�]n�I����0���GD������� �� �U(���y�w������Ⱦ!���YB��ȵ�� <"�鎖UjHJ��(��H���(��R�V@M�Y �E큋���і�v@ȁ�p�P悂�a"�+bƿ��s������^�v�վ^��.?�������������E�*�y�"�����$��/��o�E.*p�*`Q򠏛?��<�Ae_Y��}&Z�r��x�>}ް��|C�S�9�DIU?��3��5�+}��Z�DR��9��9[��I�+�l�/���:I�P$�/���\�>�Z5̝>���0��ׇh\�jy3}��W�p�ݮ��ekh��y�ї	���{F�c�~(|/DPW�6�h� ��[e�����~�1	���V�.�
����Xk�����Cq(��S���*(����W�I�xe�,_������`AKY��,��N�yy9B���C�i�k��-�1)4Ah�D�c��A�(�]-w��I�K�{�3ݨ�#�OO$j�;V�XL�AT�z�5��CͰ��ԗ��	�dTC����H�&V+�Ⱦ�P�6�s�XK�2��O&
h9�r��l�v��QlZ�>���1U)�+�s����q�q��oAT�u� ��Ah��+�!��gXt����)�+/s�e�2����<E'�u�]`�xDI����afp�m�� I!�<�>���%�ʏP�Z����[xM�"��c�Y�� s\u�Y�,I�W��; �<b*J��6*p��	(1���@�FqS��T��XSl�7�.��g�_���Ә�N�$Q`�^��X� i�목Hs�k�e���''��A︊���r8e�n>[HuU)��>һ8�g�.�p� �Q��