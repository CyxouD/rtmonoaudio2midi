BZh91AY&SY�w�� J߀Px����߰����`O�-�q�U
QI�bjyFM4i���4����6����!R    h   ѓ �`A��2`�T�D���  4     4d���`F�b0L�`� �*{M5'�	�e<� 4�= ='���=	�I ���$�'$$I F��;��_0}>5R�6�P��_&R<�$#�,ch�a"�.k�:���� tJ��1,����t�s��wآ�eDR�lcm��D"^f��Y�kL��$V�H�$����r��sJ�%�aڌ}�Km�D��Q$�-;�dw9H@Y]2$%���<�;OML``���E�u���j�i�A��wL.�P0]'0z�PD.�=������\Xg>H�/�!�,wD�9�c��9z�U��(�=�n�s��� ��j�E��j���|�{����(+��9@��%-\>�؛eP{�Th#��C�p��D��f�T����4��@kb�f�E\�y�ɺB�b]L��4���u�6��ݟ �c�m3b�͙Ug4��d�F�!�G^�g9�{�t��f�5�;����:`3�:�{2e����ec����tӒ��p@��/p٬&&Dε��gIN�j�����<�R����f�'H�S��R�0)Y��X�g��х��\41����2�F�D�!)blD��b� iv����Gn�X��asU�����$�,������~D�E9�Ũ�[#��F8J��^^{�+{�wzQi���2{-2鿑\�zyyg���	�|	��k���a�5%/WѸט�z*���[^!�%v�����<������57���.4L�����Y�z��8�8s��żHqw�|���Ϡu3j-F�H��J��F)˂K镜)A;UQ�߁U.>2Q�G�윆�����Ha%h�#k�#�	�kt�R
p��u�E����8�l�3;�{׽������ޓ�/V*ϸ����B矕��n���@�e@u��\�ڧ������zY�$��#al�I�!�-��NKM�5W3�q�cc�{Ϟ�}�"o��������,�HC>�w���3�kgM�c��@�|���i$V�P�-��I
'a74!/a�*���"�2�)�3�����Ek���h��&��n��X A
�=��{x�r#X6��Y,1
!O$�����!�F��dOAI[��5�����5����8�͊�1���Ǡԙ/��r�����|��ԍ�h3g��*�*���2�A��R��7���ʹ�[�0�m�Vݺ��Ě�%b�K�\�Xn�C�0W�UÍ�*�a�%R��b�<n�5l��:RI���D�mioU,�H!Z졜��f+��RX�k/���0�#�Z����sَW9"�L��P핅�w$S�	�{� 