BZh91AY&SY��3� �_�Px����߰����P�w@C��f��LM4�0eM3$�?I��j4����j��*h&&� `L�  "�M4��hh4F�  "�L�Dɂi�L�ɓ#MA�#A"E=4�{T�0��SM z�#!�1��� ��� �"�@�B@@���Uܐ���6+̫�HI�a@�2q�HT0D�mA�N�6,x�*B\2�xz$��:��z��/+d�������"�)����ܲ!��?��?��t�樑���1����8$e�7N�i��_ƃ
!ސ�I�� B�-���z���UM!&�~��k��{s�z?���Pq�28�mp]�
����]������	R3��M�j��/�1�yVl�l�f�"��yʛ�`:�D* ���`n�Xk�R�J�j՚��]��D�YF�B��eY����+�+\0�
�J�C�����A���p��\d��ˑ.�G*5:DC�[�!��Eg�+dh(�і���%��!.�C	��D;�p�e�$.l4�S�;�����z`��V�t�ThL|�j�'0Q����<�llm��l$��o����J^r�i��]���E������Iv�1�ǹ�T��Q�Բ aL��������,iA���a��SV�7Y�bBm-mk`m�&��yDqkh$�t���̀7ǻ��^^�̀-7�6}*�lŝ`�HK�����f*��$�UDL�$O�97�>3Օ�m���:�ғ+f�I^�ӷ/xw��`� ��=��%�Ap[�;�n��I*|�-]&��BS��ӊ�˵�O�BT|���5X9Z�����$O�Q]<m�ZD`�u.]���%��vt�&rZj�6v�nb�����x�9��]&)d� QbZR:�rk�+���4qM����e�;��r1�-W�Ah�Q_lЊo1Q=�ԨS/�ZBUv;�G��x2�R����x��
dTɏ0^LIu�KEe �/�TF��g�&5����#b�G-�Zi�����t^��@>��G'w�j���+MZ�!�� ؐ�v���F�{�7�a���,!�ǈ�+Z*���Y���Nl&�э���cR����Y#!jT���*��n�Y������!�UOO>RdgHKJB[w ߯9h����`�vz�Xv�sxB��t �]݀�t+�F��6t\�Y��$��ԄlL��k���HJ
m��s��F�*3ur�=j�jv����^��Ó1)��A�~6J����%��&3���%m)�X�OB���ny�HJ֐�0�nf�\��
Va�+��[Cko��V��� Ē'�z��X���r��<-�Qj�d�4�l� ��YF��iSP���ųt �������pU�rE8P���3�