BZh91AY&SY_$�I L߀Px����������PM�'Ē���W	$##I���<�M�f�zCj4h�A��aP� h &�   $Di�Fjh�m4i��L�`LM&L�LM2100	!�O!O��Қdڍ2 hh x%^�D�,$@�D��ĝ�<;��H��e,��IC̾�:��KGi��\�V=y,�$o�ݻ,�f������·.�ay��m�=w��k����[d���3=�b��A#3bI��&kU����P�	�dP��]��xz��f�Hlm�����������\�����r��l�D5c�ج���=K���qDJ����Z!��A���죋a9�3�QY�ɛE�`�33{	��D��Y�R%�hE�A�Z�"+@dKhT  s	&�2���� �J�d:e���I�9�,C�u�8Ao�|XF�llm��m�o.ꞂR��媽+<�d�\Ej�x��Y[R�
L�Lc��Sd��]$1yd1���_<,�.�I������ƻ���Q(�_>m�x�����+���oכ�V��D�D�ʼ�5ĳ��
I#�����Wm�-�'2�;�(٫�mdSac֙��9���r��-Kk�pB�!�w�;H^d\8ZI�7�X�&����[zQT����v�x�k#��[G���Ji.đ�r���@��ԣC�(�'����irߒ���wOH����db�Ԭ���^Y�&�@7njw���k �DA�-)�+�L)�$uߒ��L��08�+%$9ĵ��L]Y-��jF�|ٜ��qYMu*T�$VQ��6jD;bC�U:3���!���t*t`>r\&K=��tf�Vh��o1A�e�8m�"<K%Z2�y�E񱱏,^����#_V�,�k�J��fv$RGW�t�|���z�`����TA��)$N�A����84�N�0`���ri$E el�' �|#z�EEwSy��$ �(�m��r��@;ODA6v"���H��E&;Ţ��OU�����#��ק��5�sav��5��#��<��bUE�$<,�ޙc;������|���Xe�џUW�`rI\0� p�>�$(@��>Quj����n���P*���]U\����ғuw�*I��M�d�����Q��p�R��������Bs" ĒE6��y��\���A�&%9T���Lqp{��Gi�QS'�̈́[9��i��t�	�rE8P�_$�I