BZh91AY&SYr?� �_�Px����߰����`Ϗ=���` ��cA*�H&@��<�i#51�4���%@4�ɠ �@ ��� �d     ��J�р	�h�0@�2b`b0#L1&L0H�H��iF��g�L��M��Dz�C �LOR�,P$߂BA& ��'$����g�|�>?���� jR� s��E��G&�,�S]�/O�w���U��Ig��̅�t4��k(�	W��y�0�c4YQ6�c�$�jM�1!,&�^
���lqwQ7���LB��(�AÒ!��*&s\|�B��T$e�Lq�p�x$c�m3&�el��������D �۬:���9�jL��5~�a�aѶ~��y16z�f��\q"9��0�jZ��ei�SVy*�B�b+I�@FA4|������+mOhǨ74�"�$��^A3p��49�M�.$�	k�9E�����lh%�3
Ga��#�"�)�G�x1�\��([v�eP���)L��И~
;1���ݽ�5	�ƭ�5�1��i�ɪ���������F�qՙ$u��Bb�m"�6��AG�#��ZL�NV��ȕCv�i��]�k#1m)Ӌ��!���F&U��᭩9x6n��XYΤ��a)<�0u>:���iz0&Y�o(����j�S֪��Xs4���@'�F�Fr-ޱ^z���9)UIP��l8��2���+��;�c��uʍe�X����TN&���x�UT�E��f�x{{{y�P0���j��vB㾈�i�v�"��fO���壡(>�1!��jM!��1�{­�b�Ȏ�dL�^)�sz�`���n�y7/2�e�B�vE���FJ�sOo�L\�[������5WMUP`�G
��e�75�����Fü�f��fj@�b�&D!D�	��1�
�բ�R����!{F�;��Z�K��G�\��! �%[Vōv�{�.�r����i=k�GoO�О=�%�_Ǜ�����Ʃ
�5e��2�J�*A7����}���B0�T:�`Q�A~?.�5��i�yi���-f/BfY���:���B�A���Bd n��Oa��v�����Nx�,��,��e�űF/Ҁ�'� �z]�c`�-d���9�\B�hYmiD`{�+�S9۷	N	ܖJO}*���r̖w>,����'M�� k�R�e 	����T�����[v�r*1�B���sL�Y���w �c-n���e�_Z����A���Pp�I��Dan�Y Є���Hu(R�:/T_�@nm:fKEd�s��R_�h,�dO@̞��҄�Y���]�HA\|�lc�/���ʤN�g�W��<V�%�� � �w.@g��1;��a����CA��aEBw1��FE�:� D	���"(*jR�?F�H�-J�S��AM���f��P!����&����f �A�Ҥ��^s �����Xn�������V�a�yZGA�������@����0�p��Pl��C�;?d������f�!۩fc(O&�h@o#��T�3�6
��a�DT���lT-��3	(5Ykh��[ �̩Ry�����8d:[rW:B��׎�Ǆ�r[$Q`����l�@��uL�Z����#��z/���BY���FLO���==#L����_�w$S�	 s��