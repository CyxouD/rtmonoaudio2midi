BZh91AY&SY�a� D_�Px����߰����P���z�s�{tuD���I450S�b����Q���j@d�5=b������CM� d���PQ��m#�4h�� �@"���z��4�H@@ �"@��E=2&���2i����@����e�F��
�X�@���_��;{�vTe�U$���N�N ?Ef@%PD&��PÆ���e����d,���mK+����f�wmJJ���STUR�r�I�K�j���B���E#Ui҄�i�Y2Df�'��8�������"�ǒa~���
�U"�c�����'̹V��8zP��`봦&G��f�Z׊
�w��o�|8t�6n�%��� �PF\8��'<�YF4B�'
E֛��M�{�"J.	�˫F��L�M)��K�����!���T[0�d�T)�ЛzP�I7N�$��EKX
�g���tX8r�)�6rU!��b��UP c(�j$^)b���f/"��#V���4*�!̈́TĂ����/>�!�I		/"I$� C7���&#�_~ъ��n�nn֎|�<����"�r�Tg[`��k	E�Hb�aC9�ݳB��Ʌ�S�<�����P��;t%��i�,�W��-����_��O������t�F��x+�}D�83($�Ν=߂j� L4�)�h�y�Iק����Q�7!���b��a�N��g���-���B�rn���N(zP⤉��9u�G��Tr�}��b� <a�$�U����"�n*K�R�1�8��JIC�[��q�	]5p��+�j3r[;����:��C=�b���������AB���Ι[ �l��F�!٘�ңRI!����3�[�δ�A��[/M"I��B�/US_�t�/)�|(����j��L���A�N�q�R���#Ue������ �ٓ91A���#3�Rš�;�L�g����p	$R�,lc�'�7��(D��m���1�uS����̒F��VŸ
܋]ƽ��`? :"�4�I��*���i��u%{�	�t�B&(�RN�P�/�j�(�PD�	UD���n* '(�����u�V�)$Z�F��T.�T'�����(N _��J$�V�5���3���1�G���\�A
�Y;Ș%��p"�Q�>�"���Kmm�L��Ҡ5�O���hŨgz���6۬�$6�Q�lfwb��f#Ue�|7L�N+�=vI"��EsJp��z���A�s*��-ׅ�3[��Ⱥ�A` 6H����5B��y���S3�h�)%*U"΃.WT�h��,˾}�	6m�H�i�w��m�w$S�	Fi�