BZh91AY&SYtM28 W߀Px����߰����`_�u���T
$�OS�b����x&�mA���zA����4       0&&�	�&L�&	�����D�h4ɠ  �  4����&L�20�&�db``$
bi����4�zjd�S�4�4Ѡi�a��G��1"i J/H���|�z�@A��|*��0l@5<�����LHFU����EX\�gR�rц` ����1��Z8�q�k��4!(,�i��E�ў{:"B�!UUN���b�d2�"2�!J&�/�9���#I=���
�-��Gj�u!��#�0�g���A�C��!Zj���B�@e�۸��4� f8h���;3����4��}�=�=3�R|o,\��o.��3Z�mԧbN��Aꤧ&�D"�H�8էv�,���!��K�*��b1�S&�EZR�ք��IU`J�n4�,�;D���)st�r:&�܌������K�hg��֐P�jk-5L�K&A��B��2J2�2#^��ㆌ�j٫�B2���c�E^I�%".�KzZ�#Bf��t��r�ZK�*�@�$E��Kn���*ھ�y����H+��k�tf���tR�cqq�ÔVV�� ���b�;��/O�Y�TzU��ŗ��\� 	�$�ԫ߽K�$�7���:K�"��=1�,�X�#��C
D�0�K6�"#(�������Pz�ݳ��&5O�K[ZB�T�S_�}���r���lr�\��{ЗG�O������n��EӅ_Jo��3�5J` �^���yE�x���=�-��#�'�lHJ`����h6y\.�(r�~܃���>�/b.���A�!p���4��5,W��|��'\���$l2���"���"�������fmEQ�I�)'��)�$A�)��Y�o���'�T�\UOɞ��axE��׶zY�8F֔�&"�
 ��$9��N	����+�8�y��H,��Й��ݦ����c+�wDI7���������4���DEi�֘4%%�H6)܎�U��n�}��׉p/V���G8�zf�iSp��@p�2Y�6٪��)��61����X=�;�Ɖ�c�&/@5j+d�� A�δ��9�g�gk�r�L1P:"�4ɢ�*���i��u%{Bj^�s0B�$���E�MY��)�"A��L�콅D!P#�}�=��Q�@Aפ�U�.��KT�q��:C�g_�� ����WF1�=K$bcU�J0�+��L��uq � �=5�N^E���wl�JX�e�@Q��G\	�"`�g���=���1�vG�j�p���ċ�\���7�&T�~oe�A{s%4�^����R�c�U�͍׆�����uĂ�@q&�\��H����&s�J���>{�欮�l�n��M���lT�.��Wc3�El�#����
?��H�
��G 