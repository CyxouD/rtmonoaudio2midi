BZh91AY&SY�F �߀Px����߰����`��p �
�PJ�	$$ڛJzh#&�!�Q�h�d�M2z�dڃS�4%R    h   ѓ �`A��2`�U?ɕHd ��4M�� ѓ �`A��2`�D�5`T��<~��<�i�4ѣ�@���"B�	HH�B���%#޿�@����M�`�"���Rq�L@� �ch��EX`�v���& �9IS��3��n|���s��S��F�VTm#vh�SA�e������i(�N	�Eђ�t�6Jr��2h!	L�@BQF�~�P��6g��l1@�3�c�W
��C2&e%�xY�]�f
��@)�^x�"B� �sgi�)� 3]��d��kҹ4�ո�,� ]Mk'���n-#�	�9k��3��r��@��ǵ�1�dh8���U`��p�F��`X9��L�.*ф�nFU�^�|$ O!�9N��WM�E`y#�=,�XM�X��͢n%ۦ��f��S[�!����Mt����l���ȸi��ત*;�GH$�O/us\�f�f�a���:1b�Iݭ��5A��f��P�~�Yv�병�;}1r:B�l"�-�ɜ~�'��%�8aQ�ڈ���2�)ǉ��_L����3,j�L
;@��5^v�&�(m�p�N�2�oE6�#x,]5�F"�+&��nTJҪ5X�m�LqY�ڙ��,(6Dfʒ�h/q.�W�<Ä�d�eL���8��E��ͫy6	d��P�e6l�f*ɔ�ƥM
f����&�
+*J��]��x��cA���P��v��L��:�v�G�ʼ�j�<�|�ةk���fם�B�YU5���k<ݴ���anl>�_?���sm��� A�����$����Ebu
Ϻ"̓;�JV�Հ]�u��	�� !�"���� �`@\�T�77laead���ig�&$�-_{�Q����Q���\��k�ѻ<�|x�1�n��������r�^4^y�r�7r�� �����V$��R!U'�Mϟۮa�M"OVQ�w<�p3�0��մ6ſA�r�E���f�93��`��Sh�R�y%w�9��9p���Ѵt��ӓ:�Fò���� �0���8f�Z����)�OZ�M��{����u����<�}�Lp���v��NMB�oe53�8!�з������$:R�2�	�APtȎ��nb�J�H�R��&g�o:�A��W'�ȒoA��K�����r�y�.(�����ؘ4 �8'*E�1+���sa!� ��Ȉ/\�5�wL���8��\fK��uSA�4�0�0ս��A�L9�z4MDv1e��/<5��� A���޽�k�of8���0�>�tE�h6tFT%�4ƋH�ө+�R��9!�0RN��GU.,՜QJҚ�$J�$·e�TB �@��v��f4�P ��:� �ߨ�)��Z&�� 鉛k�'��5nsc����9H�9M&�jaF0 �-z��3��@_�<+*����c�ͷ�2-	e�:�e p�/�!0: �Q��c�sFȰKi;����	�̤aZ�V]WT�p�2�M�{l�q%4��gFvB��1ʬ���pӶ��0��Xb	)��?
��A+]�3�Y�W=J*���N<`?� b6�q�R�����M��	2E���(���"�(H Ɂ# 