BZh91AY&SY�� U߀Px���������PM�n;�-X���	$$�L�h&�ЙM���4�&CFM14 �!Q�����C&FF@� 4	&B��)�4��5 �@� ���A�ɓ&F�L�LE ��Q�Q�PxQ��� �`��J�̠XH���D����N�;W���\��`�#z�0��).�$��(�ѽ�EY��V�Of�-�O*�g4�v�]ڝ�9%�U �У���.�٫�\���9�F��Hˌ���{��H�r �JFh,���7gI�1Iqz�i��Z��f�>�l�y�Z�ҟ��jt0t�i�&��ԓ����ӒjMZ��-{ f@��X�f�����Fdpx1|�ظ���{���<PRK6���VeÚ�2a��s�"����D���xyIE��t�|R3&%�KQ�af4L�ʗl-\d)�a�a�d4�>��������l�]�Jy�)ty�.V)P�9b,�f�6����p�n ���9s���6�LYix�\�A�H-�,XTaf��1f�$6,�3�~P�ھ�ս�2�ش��������b(�x�>\�~;�<��|����m�N�� ]�h���.�X�;��zx;�nӏ|��\���E=E×��V�8�!cX��.W��ݡ�9|E�d6�uC`7��'����{V��,=J$�p��=�G��]�W��L��_D
=�r1���2tQk�&�O[��B� �e�K�9�8	J	�)�_8,��r�Ajj�%�C�54���4��VB�OZQ��h��DG=�*�#���A1�sR�9�W��3F��סC\wpD��)|ʊK�z��>0�����C�j��0bb����AeSN��2+�2���C�I�qPH���H,�q�͌5[����j��5Xfj��\@��|��&�.f-�B���6�.}�p��ɉ���(��ȱ�Ej*�i��2(�I��	���"DP\^�8t�8�H�W�+8�M����j�iu^r��0��J�yp�1F�$V�93�*-�&�?�TD�<�=nsY^�F`ذ�F!��k:tTd	��P#Za��q�Sj
��@���'���Fʮ�V�uZWCdU5ɥ�Y�B@ރ��pK�Qfw-��IV�n
���fR^6�jB���p@��'�6��U��ha	d �-4ŨmUs�	kI84H�H�V���i�@�
�U�r��F�%;���6g\+���2)�Ļ��{1��H�ɒ-�v����]��BCT8g�