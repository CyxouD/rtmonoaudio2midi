BZh91AY&SYO� f_�Px����߰����P��M�8�l�4	$ �h���yS��2{J=L��4i���&IP �     B(Ҧ�Sd zC@  L����a2dɑ��4�# C �!&ji�mM���COPoT&���@�	W��!+�0��$�I��̐.O��5l���j0�`M��� T`��70�����c�i˹[����,�� [�����=���R��b�A�$�e9uwj\��Jvf��%��G#t���e�*&3T�hc��
렐ʲ�s+U,3F��g!!)�� QeP�f�q��jilv�|��y��yN/�7sM��jlf8l�t�f�|���u03QㆾDb�܍y ��	m�0f*_0������*�-*!�A���C�I��h�U,�vf�.ѥ�1���g�%B�H7�Τxba�c����c��X�Zb�"��`HgH�YfJ�m� ���5F	LV�>����O5 ;$�1��b��؁H�Xoq1m#��E�� �ݜ�4�!4�/�lb(kB]�����<���	�9%���!Y��y�K���d�yWjL�L�L�`�h� ��&�aC�_&��j�IR'$5T��4�2Z����\[L00Ѩ��`�HfA[*�ƻ��)˙9UW߫E��헏�D'���t�����ߧ�s�*t<츳�X�����_O�\4��V	.�gM�9v�eBC�s<�}��Q������-���� �����V������a=F��ط����,��ދ_x����TO>�2_���@}g�H�����0�-d�#k�#�O]����k��3���%8'q�R{�'�5�m�b��騇�~��4��`�4��ĥ"9 �4�KdVpOl�Q�.?��$�3�(�jb�Iv��-�W������UJ�A};�I��X���q��jLOzpp�P�7Qz��a�j!�4��������&#��=�@|y_u�	����1�I�?���Љ]͍+o��9���<)��1�-�oB5��W��0�|`��4J-Y[����6�O2�`�{q��2Z*N=�.�I�h�<I�ĥ	a
�Jf��񙀅A;|;5��H��e�I-�EЯ|C���N������*� ���l.��T�#�r9���aN2@�
��gۼ.� NQ����XYQ�ٌjYҬ8�f�pf�N�E�"�sZym0��Ӊ60�c�)�RV>1��J��u!1��s5	��
�����UD`�R�A�s,Xa�ۂW1��k�Nc�I82 �E�_r^�Ŗ��\53�c�݄�ST��l���!ffG�z���M:��ps�5�d�lw+���]��B@?��