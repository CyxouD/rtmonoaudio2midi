BZh91AY&SY��� �_�Px����߰����`� wOy��B��H�dLI��&&�I�������aShT�      T��?Q��11����404�I��@hѦ�@ ���ѓ �`A��2`�$P)��iM�ҟ�2���)�==L�����&��QD�
`
��)�bׁ�?��*���p���*�j�s��T�@L�"v@��P4�N���ëȪ�j^�Fdci�fHMR��)��;(�3���W.K�dJ[v�5	Jn�![�S*���ۈ}i/l*�����\������6$0.�a
S؂�M� @��$�azZ����(�$��6�Krˑ��:�^�^���n�� ۾{w<��\]���x�?*���e)@�����m�!4������@2�9l?�d�D�wV�84ŭ7���4���$������v]�]�����T�����m�CԨb��kMA1H����PmC�f�ɉQ3��Cu��QK�QW��$[�ْАub�f�[���0�ț;�����(m$暠�!`T���Id��%X[��ڻv��#0@k"�V�0�!U\JU��ضDr��p���
qd�icy�e�C��spT���]�da����& ����ϫ���rBBI�I @��˯s}ů�����	{)P�#�)�����D H"��,��1���H8�u��A쁉���+?%��4�=����Ew���6w�f�� �)vb��P�i�3(A_�GϺ�~9&��D{�Bq�+��I����/�v2 C�B�ğ�d�w���<�h.��������w���=�΍��Ojf�$U����f��~��=O
M)~	�CK��h����_��ڀ�l�RI>	w��,��'�`�-b���"A�=�S;��%H���!
���/�ƅ��ɓ����{��F�TP̀&ح��ql#1�K7�\ X;�Ĵ��C�H��b�ƥ��ڂ�'o���fĴ��SQ^�)$%��ݒ(����<�V K���u� �oy2ˍˏ�"7n�>4%�※��5h+�̑�b�����9���I ��fl�m��H7���|��m<X�Ea ����2I ��^ `���V���.� �O@LS2�L\K�F3���{�(c~|���ѶPC�݊�ã���[��.Yv^M\>���d %8�su����lN%P�U�&h}{x��ݺA���Ը<�o�}
.f�������ִE<�'��;���*�۫�	���>���ZI��;i�2�����+W2Wm!&�>�;��������l�4��V���e8HU.!·�)E�;�.&uW�bIY$�xB.���0�^4I�0��m����  �ĊD��p?�q�"h�u��t��N�7JO7	��A߀k$O��8�>\[nC��M��n�W^���rE8P����