BZh91AY&SY���� �߀px����߰����`�z���@^�ر�Uz��B��&�~L��)�M20&��d�4f������@  A�   4ēE  h�     MI��4z����z� �y@s F	�0M`�L$H!�ș��M�OM �@#L#&YTGw0�H� X��G�|&� No��	rb��6�2��b]P/�Є�0EX�80��V��ܼ}6�H�i�V����Z��߯[M�&�,�T�K���d	��G6h��[K.,'��֥��?)�dh-ekփ����"��HB	��0k���ݲ)�@������=����|�Q��0�S�`�&�)�R	D��R��4���D̆ĢZ!9Fd�&	.������h_T#j���U�]u/R����c�Z1o�A4�R\P]��c�L/�E߳��)\ق-Z��
M�� Pjx"���j� �Z��m3jV���)�	0�e�]�J�c�[\`ie�B[&�&���a�)����t\*�,�i�2��5C+�q.�Q��!2�gEe�[r�T�a���f�M�v��	�$�;!qf��.�T�kW���Al�o�/i����ur�ֹd�E�6{�G3'e�0��ْ�r�%�."�㜤FLAO%�2P��"��E���3k.#\\8\Komn���Y�ޡv�G�CبM�>��K����n[ٷ���z=F�EҪ� BQAٻ��8�n��Ef�U+dl%J
�H-�H(
-U#e7T�M̓��\rԔ2LX"*���aE���b���S�,��̒CP�-g{�#/Ig��vJ���^��<��Hxn�����|;�+8(��c�VQ�l�) ]�h���'�����#,&W�R�\�~�11��ݏ�t����f�TN�����&/(��d�;LHm(�\<�jM��j�Z �z���\G����kͥz]����){E�fb�F�S'Iʘ3�"K���<����Or�+��s����S,�|ʜ���&X�^ʃ�~�{.��CS,�Hd0B�<iHs��-8'�C�+�7�>y�I$
%��.��8y+_j�2�xR$��X��l�T_o*H�p\�Μ{�����jF�-R[�xb�i��d����.;}Y�	�k�(s��Fْд�˪���$
��cc�=��`?քK6�Z��n�5�6$%̒��\ �����9B&@:"�-D�}�U'�i�Ȍɧq+0BP&��vd�LP�I8z�h���SW8��$�����3[�v B�@��.�|��(�$�,� ^�Tp�V(h�q�_H��5|�=-�}�]��åkiG��v�t��@���!g^��zH�-�>C�ȗ53�ۺ�ZR����*�c&��fD�y��#o���o�\��5ҁ�D����
 �m�'T�+�H4r9��0Y�6B��eUu��˦���G��84�H���X��Hi�@�L��*���*��v38 �H̎��V#��˄��rF�#EN���ܑN$ �8% 