BZh91AY&SYR�t� T߀Px����������P]�ov�æ�&�\�I"jyLL�Li�FMG�CQ���4ѣL�	�%O�=� �4  �  �&��(��ji���F�S@ ��j�   4 �  h "�@Se6��Si1C@ 2hhЂ� �@� ��!@��3�n^X����C,`�"�&���~��.ى�U�����EXZ�&���%��[�l٠�v1��[[V�,l�ӄ�L�c��eHVFI?�Tt�I�N�$Fl4�B{��ٙ"3��nC��c�$I�		��$u^���v�0	�fd�|�'ɓ��r�u��μ���-�"bu�����+�U��3j�ɗ2����Y��@�u�TΨ�������Heh�S�"d�"��"�$ф���t5e-�]\5�v]��b�%�V�"k;Ĭ�Z/14�1':�� 69� �"�8��H<���eV�N�ގc��\�$�d�������㨽�|M��Gu|��B���B�ģ%|\#D���"
43�̾��E0I�7�Ð�8�����Q�J3�ϋ���b���[㓇G��������l�*(��S��@.f����Q\-�(����#�p��}P;�r����o m�r���-@��+C�Oqo�{]�id3 �	 nK�x�{�SW*͑J��(#4�1�;�Mr�K4/Q�yPFK��)pK�Ŗ�4
�:(��X'����"a�I|�����%)��i�^���b4���^uM�C���6و����;j�6�J�J]	�H6A`:�F��B� 'J��L�qg)�zb��͞P��^V��T�g8
�w-\h�#�'Zi̘4
!iP(a0�Qr+\��Bcߘ�=�	f�Z���\a�4ˋ���b�a��>�\q_�F0
00�0���O^0m����!<����5O�I�-��0��m���đ0�z��h1�&�h�FQ�4Y��(���hA!5v� D�ED�`��udF1h�uy�*I�c�'=�6��\'(��&�U%�`Xͬ�l�EB�<�h��=e@n��{�'������_��6���f$��qө+!��_��2��+ͤ+��[.�t��J��6��	��i,�F2`H�����%0o����4S-.�s<v�:��0�D�����\�CJX�pP��R;�Y,a
N\C�X�W��D	�$I�W���ް��2g�=�H5��+�EI��Y�#��d
��Jb^V=���$Xɒ2�;m��.�p� ���