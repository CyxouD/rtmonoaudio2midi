BZh91AY&SYm�At T߀Px����߰����P9�NqF�3J��MM4�e12�Q鉤l�C�OD���$� hhh 44�  !�d��=M<�jPj@i��0L@0	�h�h`ba"�x�&%i�O)��� �24	BY�)%v$RHD$#��'�|W@w��ꙃ��PÛ��BA�`���na�65�%�э���Ejˀ�:�@S�zKgx�C�W�z@_�7dӝ�8�FRvՎ�
�`Dc�� �V�;�܂���␑)c .����N��L�0��u[������������ ��GQ�sF�4��o�r�r�QSŁ\w�]Z�і�k!f7T	 ��9�Ѐ�E�;�I��Q�(��BB��V��Z'(�Y�Y�dB�`T����k�MV���I0Q:5�GQp�U]VOm��R�- T`�~z��s��H$���l/iN�R��l�­>��Y�"�\�y,�2�5R�cA��nXD2�ӘL��a%���)|�(0��y���B���Q��wd��%\�ׯE�<�ꗿ��!g'�
����~ޞU})󞇑�S�{��_+�_�y�'u��y��y�G�Ӿ#ƍ��[g�"u|ܩ��1@�Z=�tj?��/(�46�A����'�����ar"�|O�����
�sl޽F5� >��W䗋�h�:�d�����H��Z��Y������]o}���f᜕o���'!���������ĦN)iH4�ld�W`��J���Z}�$1�
�O��jS��v���c)v�B)�KI�U5�u�T�(qw��D[>��`�)��Hi��)��u|�]��!�$���HN�2&`BG����f�� >�=z���pa�a�{m=t�vDs���Fr�cu�<,52H9 ]�P9[�3�ng�G�9"�4�d���cE"C2s#�BS��|�,b�8{�l���T�qe�INI��n�Y�x/1q�`�]u�m��/F���h8㠸P�w�>߇���G/��OAk5�scn�:��r;�s�zT�	�R�2.�Y{�����gsT���=�[7�k�P��I÷j��A�j:�p�n$�n2���}�f��2��κ�R\��P����qsX�R�����b�/
��[+l�d:R��� �U���ꋛ���/^3g �͑VeZ���9�N( T��kQ��~�1{1��$bɒ6��W���w$S�	ل@