BZh91AY&SY��e Q߀Px����߰����P��f�'qFƌ�T�$��SB6�&	6S#OS�=G�I��ɐjm RS@2   �  H�HJ~�z�  � @ i�9�&& &#4���d�#�L#S&����4zOP  ##�
����;	$�$$���$�'q������Ff��F@	�a_~A6~�I+��Gkiak]ˢ�@L�{3�Ei�V���sfqU79L�1URH]��˪m���?��k��e�mp��?�
렐��4��}�+aڃ �I��%</<I"�m�2�Ӹ�I�00[��E���Z�:ŉ4*A�c�3e2��ٝ�y�H�ӭ0Q~n���k�5fZ�(ׅ��r���B�^R�h:j%N�V?�,wku2��'@�l�FD�wجL��2)��eN+� �.���2�R(:��]��{��xKV�iM� ��b��cPsj錴u,�M�-K��Qe����}���3� KQI����XU�i�Dh;=Ӷ��`=o��*�����P�����<����"'���`�
�&^��r%��vp��N�VL��U�!��I��I��pc���M�P�7�C �"�	��
�A��ٌ+�X�I�>%�,d����-S_��Ҏ�Q����+�}WLN�^�V��xy{>X�<7�%e=�^y�%Znr) .������)�b�ݹ1?|�5�ò�:��d�q���Zb�̀ZW&�x��?�.�1hlq����`�����йo"t�؜���U�5Ec���E���c�ew>�
[��cJƁy���g�C��]��)r�Kvs�l����F/}�V�v{^s�/R]��3��k��FF-��:��4�Kd_8'�A��o30(5F����u�LϘ��μb1+w�TI7���ٕT���S-�oq$���T����4�����ا�L6�$�R���@���\,�9�OC`�Y��&JfE��s� T�K��~��B%���]om�g��r��[ �}x@����v=�P���DXCA�Iڲp6�4e
�ZyF��	���|�,ah�t⤺�H�-��aL��H �TI����Q �P#wm��?{$r + mdP{��+��Dׯ�T��F}��OAI�C�˯h�u�-#Q���u+$� �=� �t����s��ր'.���;<�[]'V-�`J��h
1�ݫq:L���M��KwZ���̣,���Ju�id�Dy9���d@f ��3tQ��Dgd)XA��Ug�}��̙������A`D�+�����[�ɚg���܃-�I9^-���d����b\0c{f���v�GFp�.���"�(Hvh��