BZh91AY&SY_�)� �߀Px����߰����` �p�D
��$�5=����M5���LOD�4ѓ�ɐj��&�Th4� ��M�挘� ���F	� �"����i�H@ �  � hɉ�	���0 �`�0�""hHj`O#MLS#�F��Q��!O��$A$���@��ģ���� ��~w)e�6�MCA,�y�HK�.ch����V��z��u�^�[n�Y�A�������q��D�MZ���L�\C!�	�Pd��_0�I H �,6.P���1�r����)�$�yIɪ3���=,0�Fc��4+&Y+Y�ʂ��=���@���L����f�2L00f���L��K%���&�� n���ٚ�#�� :�]��]�bwI��Be��Zl�"�e)�6#�mR�bC�".�.|'�x�Aڰw�A��wF���M���!3EWG�W5�Hk�0��jM	M�q��r�*U�S�����!fl�)��"�{N�h�@��1	5��J��xl�HC�|AB01���]�Ht�V��,��!���ջ����܂��n(Zș܁���C���.�nɬ�cGVIW1g
sb���Z���!Cr��D��Z����R���E�4�P Q�Gp�ɇrg1�Ӌ�f����uq)����kn(mՍp'D�1Bx��j���D�R�Q{�Z��%f�z�U��z��m�V�m,Hl�Aa���\�0H �D( ���S�J__�V�g|E̖w�V�ѥ��b�i`w��%�����~�Id ���P&/&3����T,�Y0�(���!��������uʞ�T�{qp_�u-���O
�	]��+�y{>X��;7Β�W�xk���� ������'~�LNc���y4p��x�F�����91�3@����_0sR̻��zډ�C`!y���_�<�����kER�ޢI�NC](�piɡ�1�@s�=�~��X�,j.Gd�W�R��g�E	ke���qx�_E�pY߰���ݟ3����k��4"bJ�GKIL���N��L�7Ap:��ʕ����5�i�oE����^=3`&Q;ʅo�
�v������<X� B{Ӄ�<2(Ihƨ�p@m��|�KD�|x3�xF���"f��CNx�`���c B�\�lc䗴�l�������������:�B�འi���x�[�E�TX��Y(�UU)��1��F��؜��xJ�߇!"(,b�8|!j���TVqU6�("B	�D�c��\ B�P���}<39��.���A㻔�T�L�j�?YT�5nv��͒�<�0kXY#�9�G�ZX�B}8��7�K�ȷ� >��Q���n�)�d͸��5jU�,���@�:�Ce�L]*��*e�"�T>1�P�����ės���+��V�|���a�%R��B妙_�rs��"���Q"���iS�9qj a���l�츢�J���u�
 Bʹ~':��Ǘ�[7�$t��;3#�П�]��BAT�p