BZh91AY&SY5�o� �_�Px����߰����`����  :��@��I!��G�Ai�SC54���� �� �S@�F�4LM  �A�ɓ&F�L�LSɪP���#L �11�4�dh`LM&L�LM2100	LB4OT�)��OS)��� d�B� �n� 'a" $	�B		  I��z�H ��������`�4����ґ�Q �0�1�pa"�5��m�ާ@����p��C67Jt杖'�76�0�
b����)�-�[2T�BA�3)�)6�pRJ
?��>x4琍MP��ٖLq��f��x�D�`����� �W"@(�i@$`/���>ߑ�I� ���O�8a�z�\����F�i,A��dŶ�D dX+�[!Ę�& aKE�1z2 �W�v�BS,
���f�N��.��ضi�;5ԉƪ����;[���a �E����c �1<�X�R�>���A��ٛX�,��M�d�,�7Ҕ��c:#�	�PRe�e a3;�i<5�ޜ"��ɋ��ݭ�)<�PN�@�R�F]Qb�K��ͅ�!mlH���7b��͵`p��:Ӻ�x%�Yj��c�s1D[A�`��лD[�vg2c�,�rXO*N��q�yJ ��@�e������0�N��sM\Sm�6�I;Z�̰�L"5�A,ћ�{��6-5%��!� �<���Ш��n��:����T3��܅ǉygYX/I:�*M� ��SD�ax�Rh��<V����u3�6��x��x��̖/ĩߣ��z��"�g~r`Y�׹�<����a`��n�N��5�(�l۫��5ET��uqS_ϛ��񏀒	���I 0@A6xt)�%/���Um+=�2Y�Z�z0���{I" ln��!Idd�����b� /X�����-\�x�Y�����3��7[��4�ݎ�C޶Ǫ��rMF�+����~{�g,8��Qk͛�<;0گH �h�����4r� ��I��|,+�W�$�ƚ����>'�F&c( �|Zd[���+����@���.�"x����r�D��;�C#���6Ic���Yt�����?��H �Z]�~��4Ō�fzD�D����{��_>s�n�����*�q�dw��$ �NCO�X���[W &�A�Z�&jAM�X������Tj�)H s�g>tŔ�X��A`���3����I�N���� /+�>�G�$o��g2`� L����Z���=�{��ql�Һ�@�ݿ���!
�I��2|��e	�i����P�\41��L���P?
�7��\�{Y�n)�$;���؁Ԁ>�޸��̲=���@�}@�Hh9��U'P�-�<t�Nҙ�S�]���/R�=Ѝ�H�W*+\U[��b�g3�q, B�GWA>��M(�H ʐ��E�1�
�W����*��GS�'���1^��aعZF���;��b��i ^����p.�����U�l<��u��Ͳ�����,��T���LJT"��G��_f�rL_*θ(�<�eAP�O=j+M
kh�,:o�ؐsH �$��zΌ�6�d4	ՖU*ۨ��)���A"zƾԽUkO$-]T��h�1�E���8; ̎��4X�vL�q��2d���Ч�.�p� k��