BZh91AY&SY�� �߀Px����߰����P��n�!��-U�(BI�Ҟ���ښh52M��4h�j��3Pj��h&R� h 4    	��eL��&���hѴ�xS�h8ɓ&# &L �# C �$�R��~T�R{TǑ�=A�F@ %	,���$�ĊI	��$� I���� �W��uL��`$�0���+����`���<L!�Q����,<�l���l���tAN��ŸW-<x�Px�us�.ͩ�D�j��1��m6���M�N��*�IC8+]X��ٲ	�456Q�+�� �.�r����H�,����'GI��`��Ƭq�<��ք�����_j�ᱜ�3e�2 ��%�Â�u\+��"0&��(�JͼL�Ȅ���5��9�Lw�f������"��N<ު��X�t.h���q���;36ף"���.�m*&U�1�"���wݬa7�!,��ԇ��5�P,jq;���V��*V� -3�s,Ywj�QNI��K��N5��T �8D�M��ֳ��acR4ZG
�ld���6c���64(���[1S'�;7&ݲur���s��66���m�@�M���?�)z����V���Y�#+�B}mK���ɩ3+�a�#J"b��� �K����yjk6dռ��0�3 ��mcg�wl弜�����>t�xf���_�����~������������׭L��q����J�Ё&*���`Q�A^��|G��޲��̾�S-fo�Kya�ܡ�G�� �Ɔ�K���廰Ma���s-")G���!���Y�4y���ŭc���*{�m���梾D�*�(�'��V��3�a5���v�D��JO}!d����2�����!���{j������
 �KJA�V�M�p�pv�3aϡa�4����arb�In.W��\3��.zf�TQeu))�ǌ�'�3�R�TDW�x�R�����>hʌb�I�����`�i��*4���L�s�2���M1�}�� ��;�lc�O3����������nV&Y�*0d����] i�j}��[�"��|@��^HT����m�hđ�I���SˍI@2�JS�g4#�d���Rx���INI��kQ&`輥b�L#]�ɠ�m�р	bZ�� ����C(W��{S�:�l��
� ���6;���feK$i��fII�0	65lB6��&���	9r��(H��Ok5a�jY��b������%g�⩄g)�����گ�5�`�T�>PR�Q%c�ؤ��:�	�(5�kPS`�v`E�v(���!ţ@�]us�3�MM�:sI��A"��Η��2� h�p���A��E�)�f5jpwAV3#�`�&'�~2l�H�i�eln�,���"�(Hf?ƀ