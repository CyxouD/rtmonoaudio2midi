BZh91AY&SYT�Ѱ L߀Px����߰����P�96pGqFڡ�W-	$# &��	��̄cH�� ��
T���h��  �� S"F�J�ḍ@�14���s F	�0M`�L$HM	�z��&�I�A<�=##ЅN��!N�DI� �BNo�������Q��l`jxT�@��J�,ch��E�-k�г���Kf��(�1�*���Wè�q��j��Z�%�j\��؛�%�T�LK��GF�%=rv�Q#+f1��¾�$2�L�%14X�u����$�(���4������|�Z�l}�xS�7A�»^��I�V���/V�����U�!4e13��a�<���q�nٞ�P�d"t�Q������ӝ�Q�S��&��8���Vd�U$K���6�R���:=��*�B����#"9xA�4$�Ҕ��)3f�&.�T��3�yEW�E�G��(L&P�9�ŧ9j8�J�E(�����lR��e�HVԅv(�`�Ɛ�3I�tI�Y7����z�i!!%�I$�(��sv'a1�F�F5i�oJ8����>��i����D1HH�(����u L[�P���q���SZ��d��fH��b��k�%��M<�0��|����a,��*�����E�~����u}h��&�*t) -�����)��1M#�(�>�ɵ{?۶N@i�+��v��_������t�\]��e�ú������������B�r�Vjm:�;Q��S�7���5�#���Yx��M)p�(�KS���:3�"k����e)��n�9�:���*����X�=�0F��8����Ll�����"d�*"A�J]#D���f�u���HD�,���
�-[�Z0�j��L�
I�N����
❁�R3�<��^\��R��Aj�s*\��ȧ�x@nLd9�KD�jǋ9H�CAa�&3����S%��&T�r�
�8X�ǔ������պ�۽��jkL�㍤�� ^����G:o<�[�"ax��*CA�$Vjd�cE�#i�Jք�	�w�B&(Z��s87�dE�bݣ0�@���ic�� �P#_���&��� \�WQTz����L�����A����J� ���k����ڭiD#��v祊ٱ�'ͣj�2N�vи��?_�č�R]�&���X��8�X&���F|zI�#:<�ng4�iv�Xa�n'|�N���]լʮ'���B��ձ�� b� c:�΄&���6!0�j�m��{~��M���@m&�f����t�&p� ���{��F�%C���>w� ���2��Ļ�f{1��H�i�k�7����H�

�:6 