BZh91AY&SY�� �_�Px���������`~<}��9��ηiz`�I�ڧ���~���HG��A�LFC# �� �����     0`��`ѐ��&��S" ���i���Ԁ�  z�"��bj4�CF�@  4��@�4&���)�M����Кh��TJ{�$�)(*�) ���s*�\�S2�<@'�C$9� �$��I �A�PB��Q�k誆���%�0�\%���WQ��O��M�UL�*��aB)��JO�Ʌ(��mwgj�r��o����$ULIB7�V�'�8�&H�Y����v���A�\�r Ak��$�"�Rv��O�$�I ly��-��������pt�@rk|*�ڜvTe1�ԫ�(Y5,��afy�|�D�EC��.�ۊkTwdm� 	D���VC\��i,%��j�h��šB��Q�LEY��[h^�t�[��6t�4m�iXD:�-�a�ʇ}��Q�4E*=��"\J͡�I��++���-2i���æE�b�ȼ�P�Q
1�@Ub��Ir^)/K�*\<�G*����*a���2QuVkb"m`�cP�/e/@5�1JH���4dd�\.�s���1��@0��f�H���ub:+C�-�(ꤊgi�ˉ�<-eJ��o^��!!%�I$� ɿ���LG�ozхZ{����x�`C� Y��J�m&>�5��
�0�D�" Y�Q$���aU������aa��W����M��K���D��Jz(��v�S�O���v2����Y�|h�����Ys��vb�˚x2�$�vU�ϳ��]��`�L(]�q^��eIr2��͗��)�l &�f�|A�x��G�P�
������wO&�z�E)t�sD��+Y��B3W���� �q;��Oj�V�Y`�sH���d�.�EJ�g�J�ao�z��Gg�J�(�gkL೿y�F��St�Z�;�T�Κ@đ�ԲX^0�l}�$*�2gL���+g�G.�aEZR�@�"���k�n�U��#Q���M�)&��3+��T+y���BLZ���@T�@4.%#5�
�!��G�Jd�i$g�e�\_�S�3G�����m�k��I �[���\�)����	�6�D��a�?�W ��bIRH6�\�W`f�w4�|��"r��}UI���i#R��ND	���RDPT�Jp�B9j���TVqUh�P ��K7;.�����'�Ù�I$I$����ҡG<i���IRdg��d�\ �׫(�iW�E��h5橊QcI |�s���p/˜6��I �^����-ɞ&�>�q[�<�+�T���e*@oC��87��D���zS[�j��j#v�]� `���w$�^�H+������Ր����]r� ۿ_/���P�.�|6��Y�^r��V����-�c'�H�tL�7L� X�"��uU��.���l�$ci�f��t)��ܑN$40�,@