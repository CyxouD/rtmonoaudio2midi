BZh91AY&SYm5�$ �߀Px����߰����`���q 
\}檤BR����2m��5=OQ�jHh�Pɐjz*�����h�� ��2b`b0#L1&L0i�	��  h 2  4 �z�e12bbh�ɣ ���CD�S�M��j=�i��OH�����(l��C)qPZ0(Y�~/�����o�H	∄j~E���l &0�; TS����v�]�BpM��qËG-����OҘ.�vn�mZv�K�CVM�2�:�u09�BuEܐ
�LQvՐZqh[�Hi���)SCi���K�p�y�h�R��}��+�S��X��n7��۵��[��R��(�m,���h8�}��؈����{6x�^Ν�o6�k�(8m���ǌ�v�,;Y�����]0���A@�-F&y ېag��JgzN$�.e�ah�t�9Fٹe����c�4�}� O,7N:�.se<hJp�$hhT�����nU�X4X2Q�F��	�I[�TD޴:KB2&(Y�5��c5�ˢ 8��C�6�� �����c#b�R!�eyu�f'S�lO	�Y��ňRȼx,nL�ʺ�5!Źem�������k6�Ѩ�S�Tb�Æ�Py�.�C��"������f��Ƀ��f�2p�z����"�r��PM##K�8�*m$�Jѩ��d�� ����Xi�z��q�F�q�h����!��VU��:�7h��1��,%8�N��W��c�8���mUS
H��vwmX�`��X�7+�������fd��j���Y���q ďQ��;պt^զ�3h������[`ڭZe�����پ�t���N��J9��P��xů�
�u��,i;!���N��Z���~/�|ĐJ� B�P�MN<}H�%1�/ƕs�o�:���a�4t�BQ¨e�а�\B�� p�n���ؘ���^��N�3��	�@D6�Ѐ��폀� #ޢ'�,O
JD�蜐O���j*��L?j��ہo*�����8|�_R�:��9[�/�%	wq�{�@iN�ȭ�y���2�cX��������O�?�`�$I� ���p�ӛn�^��?%D"GC�ӥ(��.���jځ���DC.��!�ϼ�ƲO=��z�\�{��"ɘ 뮥ﭝ��"S�~V�L!R�}e�)���[�Ѥ��_�;�DPNh�����U�8��ɣ)��.G��J�r+=m$2Re"�Lyua��]f�'І�!���
�'��c�G��؈������^�yz<�<( �����J�p�%F[#v�#�5�XL٫N�I��Fዛ�8��)Ռ�2��C��y�i��Ü����mb�Q���P�}>����8�:�D�%�a>P�&MD98�p-��"eb�.�Ki�����,%��m�A�OF
h9�r���Y��[�,��1�'�G�0g��n8'R�$!�z��f����;�g'ШQAc6.�n�9���tx�v�S�""�oN,-(zx�@�tD)ǫ+Py|�v]Y����b���j�`�I�u��ID �q��5�O2lk���U3�B�����J�~�&��M�D3��a��^�ˣ�k
P�r�P����ꪶ�ỳR����E��)}U�aDq_�l��iM�j�FX�v�|"$ �fG�d�K�Ѳ�'��F�L���݈W���)�i�Q 