BZh91AY&SY�� �_�Px����߰����P�8�t�(�ڀH#@6�"LO$&�4�OI䞣jM5����P 2i�    "�)����H�   4�0L@0	�h�h`ba�6���6S52hz�� h� ����Un���)E�@(,�=�����\�
���Ɛ>�-���@�@K�"x�R)t�����ϓx�c����:�t]����sŔ�Ajni�ʉ��	�	&
[���qi&K��m��SNw��j�cf�8�p��	� �O0���gut�X���=���wewsz��z� ��>4�����/�J?��4�e��?^�ݐ5<i�u ApF�O���p�:
��5�L�D J)����4�3�2��a�Sժ��T�^�Sv��A�݃��h[��L���B����P�d݇)�<C�A�� ,dS�%Ui[^�����㲻$!j�<F��	O[bR	b�c*�68ռJ�D�.e��컷�}=�ily�)��)�X���g3F��h����ۆ�	�ʪ[��e�2�*9=|�O1��~��m�@�M��E>TJ^�,p�n��%�x&q{>V��rq\m()�>�l	�b�,]�18P��B��p�R���4C� ,�1S����J~D���n��;W\����Ж��
��>������~��uwQ{���S��	x[����)�2�qK��Qo	����vDxѨ��*~f��9��j@�u��s�=g@�;F��@�I ��.�-���r"��ρg+x�#�tg��V��1��]�%?z_�|l%��:2zDu��+jH��XIwhg;��%('uW<�}\�,�=���=��.�D9-��i�{���E�##<�!��`hҎ��Ʋ#%O&}D�Z��_	�ӹ�!\��T��9��&6�ׯh��Xe�X���3�ۂ`d	=���=jP�7M�M�X@n�I=,*$�����Af�D�b���@}j��6�@�Y�fk��O>`otG>�=1�^�-ʵs��C$��\w�`9�Rpn0����4�b��4Ƌ�
N��Ѐ�5>�l$E �)N��F�$f,�'��,D�"��D�}�xK�� ���o��К@]���������P�lC�����ܝ�Y��՘>�Ҥ�v�'��y��}��-�;82�"lad����ڀI�>��1��'�]&l2�*��VF�f�N�j�D�A�i۠��FD�+�+�
yePT>1�julh����c,i�JLQ��`9��*(��'�8�h+m�T�QKi)	�pm �5ci�/EZ��@�Õ,�p�a=�J�#M�͎� J�dw�Tgb_\���t9��2FU����W�.�p� U<,