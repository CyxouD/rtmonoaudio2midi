BZh91AY&SYqEZ� �߀Px����߰����`6�� �}�Uv�9��D# ��6�{DM'�mGꇤA����~�J�F��� �d�0�*y4#����@���2h���B�)� h�4�   ����24=G�= 4@  (����i�yM0�P�M�ѣ�h�lJ��ƈ��KQ(�+�Qi��?�Q���k`H	�*1����6�
��H��R)l�ź���a�b�L[Д}�ò������ᦣ,�7J�+M�V$�䔉Sr���UHQ��unM$ܹ������W������C`�e1����R�@b�d�^��n�2��rUK� �c��M���n��*1���n������N��%p|��l�(�/�z���]E���M��*������ʀ�4��2;�PF�bx�7AT�	��pyH)@�$lH_���a�k/V̪XA����Ekd�iMF�j����t@G\�xܶ7B��,1ƻ��.͆��9�"���'f��]
ӷYm�f��?fe�T��D�@�h��(#�k�Y������@T��2Y���Kʆ��Kn��Xw��nP�iz�P��4EB�Ekļ�5s92��+d���jy�I2��B ͇�,2+���c
�10�7b\{2�����ŋj-����Ll[fL��c�<L�:�Q����haC]zY�m�y�/8vފ��9"�$�a29���>��n�Bi����sl���H�zo�C�JSF<rCƹ
�+�F^sO��-9j=�_vΓ�$$$��HThP���v%W����h�_�"Q�o6Q� e%��ƄXG�����WJ��Q���J�vZ;�. _^�����q,	��A��
��p
��>#���0%Gˍyf��_3Q���xZa�N*bH_�wz|~%��$�G.r�%��	t���H�Ҽ�K��z��>|]��$-�^��]���<�xi� ��IG��3!�>y��H�T�O��#�x�_^���1�DR}"�wP�$�gRb3F�s�4X���Wї6B��A�s_~�w�1�S�0��B�	�1稝����[�fxuYB;�+
�/"�J���U�M�ev�+ރ�jv�� -DA
o,Ω�з�U���a�.��x&mEŘ_r�I~�Q�Q{WP��d��j��*���,&�c4r�5f{�#xm#�5��LM|
���D�����$0Z��)T�	!J��36Pn'�`7���:�������ʬ6�K��^k�]7����%h��\R!���o�����a���Xˊ�V����TK �#10�#���q�f*0���j�:C�h�/hU4����0Yt�4G ����Ps�k*(���/��;ì��'ؠ��l��~~}��{�M��8M�\�o�Tf�=@�)�3���oBu.vB��̷~xƊ�l������bI8�ľ�� ��p0�R�Bl��l���^BvY��r�S�)�X$�6B�l��ETU�P�s�X�[�@�:\ۇ���8r"�gG߭/�b����ֽ�3���V��STto�i����#2?#z��O��²|U���i�S�t1��ܑN$QV� 