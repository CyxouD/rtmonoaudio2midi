BZh91AY&SY'�L` K߀Px����߰����P�8��Gnj��� �@ &�dS�=1Oj��<M53D��4��� ISF��M�i��i��ѓ	L��қF��6���  @9�14L�2da0M4����"R&���m)�=Ff�i��hA��F�R�FQ�
V���mBӴ���o�Ƹc� & 4���WJmb���',
E,�lx�<��׀:*f�	G�1U�p�Z��=�LS'���-6,��Sb��ͷN]Un������6~��S�{�(�7�B��,�"����d�M��`3����YjK����f�qم� d�����>��ֶ���LM�h/nχ�=�R�ȴ��!�᳌��&sw�.s�.�u&|�(P5QE� vfA	��d1PjZϢfM�U�ꥡ�r�Z�LJ��*!	&��Y 2P$�rg3�T���4�@��^��b���;���H0GH��ؖ�EI�J����@�­Q[`n(�$[��:<BܰbCAUoH�Xz�5�l)5T9��P����)dGJ ػ_E�8�����<�SZHHIy�I$
 �2o���b<��-p�moJ7`L�r"��2�����n@�P��pJ��-� �@��C�W1�Gr6���n�z"�)�!�w�����	������|���H���<���痊UL���]�:�[�W�Py����}
��@����U_	�����F�Ǭ�,����򨽘� ů�~���}CiG�;��$�aD$�����}:�:���Nx�\��q�?�ў����ۢ�{
���+�����X�)�8��ܾ�U4^{����R	�V�o}J�b]٪���{'7�?��LA(�Q(2@�h
[D��+c.
� �dw4�E�H)̿[T#{"|K׊��}ع�QY*�RP__�TG!�4h����� �����ڡDo�JYn�bC��ca@]�ٕk�����͈p��V��o6�
6ka�a�{h��Ds�����vCV�ތ�C<Ut <�n�3Q<p��6)pPh�V��d��E�(B��;��aU��Ư�;ʄ�b-je*'���*0N�8MC�&���.@AL9��7���� � :u����1�k»:b�ޔ�;�p��Zz�݇f�0u-l��r=g	�FX6� ���p��Pu`�3�'(�I�<~��[Y�-�jJ�뢻PI�"�i͉��מ�st0�4���i�:iTX>1�Ip�0�Ly#Knl� �`+n�\ò�E����.���J��������pp �+Fۀ�p� k�ʶr8ߙ;�NF��p| �W3#�mQ��|�gc��H͓$o�w.Lkf��w$S�	�� 