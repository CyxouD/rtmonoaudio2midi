BZh91AY&SY>0�& Q_�px����߰����P�8�(G30�4��ѡ4G�FQ3J<���OI��6� j��F�  L�4da2	����S���O&��i=��i� 249�#� �&���0F&$L�Ԛ���jaF�P� �4����	!U�I$�D��I�:�t��tSeX6� MC
铈7LI+F6��!�Q��l�j��ـ�.�p�?
���?t�+�/���U2��{�,���׵+��!e�e��Q�����+F�P�r�f9�qk�(gal2��e�� �.ۉR��$��xp�o1�M�&��^��ϟ��k_��;߈̃���bO�C��s#oԺU51܆<��rƺ�rU��V��Vi����Q�>W�oE%�qlj�"�\1�E�Ђθ$A�� �KN�a�0��d����.J՘xP�V��W��}$a��K�J2�ec�U ��`�rL5�\K�����C�E���($+TfK�e��\���%�e\%�EVz��B�dwjeVr"�L]���Z!�I�ڵt��ח�6� �I��I$�
��\��R���t]bׯ�2��K�#���dM�����X�����Սf֘ M/FKh}����00ͫ�!��D!Nn,k��=䩮��5��K���~�p�^���~��o��꠸�?eW�����nR ^�����խ ��l<��xPG����Dxљ7���KOkRuZ�6���}�a�W���W�-�.�l�y9�����A)�����+��H��7r��a����S�KŌ���B7="!E4;��DJk�Eի�����xv�*���7t��x��]���og]��,�0
��;�:-8'�b�Q��~s@� '-�0�W��w|�;C\��D�x)l��k�h�]Ĵ�,��4a��P�ps�[T*G-�1���Ӊ-I�ca ]X��Vq���D�b��<�@}�U8�����0�0׽��7\G>���]lf�W<*8�$���Ҽ�\�q75gKf�r& �ET4f�K�ƊH���Ȭ�PMW^7"�2�j��Θ�{�h,ՓėX��,���px_���QaPϮ@�kѬ` ��T���ap��'�C����òG'k�+)QAa{��o��fuS$qG��rhJ�c O=��Ҡ��i��'(�P��N6�eǔkW�0璆�f�N�\��� ��o2��2Le+OD2�"����V*Uѫ*�C�굨 R`�C�V���r}#�F�B��ʠ�
�lGJC���(�loK��Zr�6B�ﭜ;r(�R��a��']�f��9U���n���)RG3M#�i�o��ܑN$�%I�