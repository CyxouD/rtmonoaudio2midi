BZh91AY&SYi�z _�Px����߰����`��;� �ª��H�S�4ЦmSd�2ji�#F#M4�ɐjy T�F�CF0��F�����ʌ� �h 2   9�&& &#4���d�#hɉ�	���0 �`�0�"@$hSaSڧ�D��~�ѓ& Si4�4�G�� ��H��	 ���!(�?5�����Z���PB�a�sp/	��d0EX�;�CH���к�:��B����L� ���I�S�޽�^k�R`sU|���ؕ*b��ZSb�MeHA���Q_Z6Ү,(�;(N�	Q4T�)R�%�ZQ,��!�p�y�e2C3��c��C����2��ѯ�a'�$$
�ĀI��:���<;.��`����+��lҵkw�4Y��n`�v�u9��vz��,��,'��KT��|�Ԓ*�!�R	2�D�8f��~�L[�D'�~j��x�(1CaA�8��By2�Te��A6���B�1��k+�	
L�h�h��_�NM�jV���	���f��y�H�۝�b�e%��5j�SF�ci�d�<��Ɩ�u���Ӎ�X$�"��1�i�1E�iN9���$OD��p�x�2�m����v�h�6�q�a�t葠�M"�l܇��q��F3�46�9�8�շ�s��h�WaI-�<JM0#e����U�ۙf.�XC[��4g8��Yl�TP�*��/!���<c9���]8�{��Ű7����6g��+�n�m��S��t5s9�	�rb�У-��^y�g��*�[�ś�\�~��߿�,��] z��*jB�.���˘K:aN���ʹ����7"�X�Z*�iqwɀ�R6ZXu�w�Q�����Y��66���lB AMHxC��˻dVH�Ro�u"H�@�`	Y���+IiC����(�~�V�m&�1�b�¦�9��gC&eO9kYI�6&�moc����R����C�@����]ی����������JV����%����e�}<|IYh$����*�^o��G�LɽqK��l�ľ�p� 1,?N+:C�-�×:/Cb n��'���:ݭK�%�1��y��S.�_጑@t����r]]X�f�Ud�M��ѧ%1�([n��#���Ӵ�>TIW{�8b}d�7���c���,�)1I�`b �#�	Ntč�}pT�#Ax�YH�R����d������r�2�{�D�z̊�U5��B6w�_G�Dq�z�&!)(�wGUw*���i>w	%�Ap]�N���y>�H�ٸ9q�)�V�o�]G B��cc�?��m΄K�-2�6uhZ�+�s@�q��}��ι����Vgs�r�L4������z*�4ƋH��ө,4��Խ��HD�eԓ�g��D�
�j�(�iMA%Uf�e�����`O�n�b<� 9wA�&�Q���=~>��tD���I�&�k��-ՔfK$c�擗5�(��@6I�iL=����*�����d.�#o2V�0��XU��G.���0oQ��:g���v:o��MZ��,	^�Ҭ�'��S"�,f��BB��d8߅��
V �s*�j�|�3{��"�$��Et���>kJ��:'�z�p����%�+�B8l8���!��?#�����f59�2d����hK�.�p� ���