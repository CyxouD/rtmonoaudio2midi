BZh91AY&SY��z �߀Px����߰����P}ޗm��^�h��$�S	4�?JbG����?Tz�SL4OSA��ѥC@44     )�	)�=F��e1S��4�G��z��MT�)� �4h 4�@  H�@M5�)�jx���=F�����43h�[��T+��FJ'�ŏ��� ;�uե@�1@3���K�����`���x0��V��̺��o� n���F�%O��K��g�hir44����4��V�$�)/���v4�/ΚHC&D'�;b��x`KAt,k]>1
���Y\�$�a8j����`�9�f�~GW�k��6����͡��^�hߺ�դ�d-��9y���'"�&hl�lX� cu������,�c��BJ�.W[U�bGċ`v /3{V�ȷ�2M��Uޥ9���\]�גE�jH�R%qCJC�	��Q�J*,�"i�M��T�Ml2'g3��P@�`N�IQh��������!!%zI$�0�E}�9؆m\��5��V}��D#M��T��"1ArgP�(cG�
LF1 �0���ݚ!`���֩�,�S@3b�����y�4���N�j��義�Bd����zL�~٪��<�Փ�Z ~ym��z嘀e���t��ԧw_����L	�\����_i�1S1�rvi� ��8�]h�46 z���_?�O��n�Z���]�(�-p�Ƿ?â�>�qԸ�sA������hS*Ld&�Ԫ��߷s%� '��<�Ds�eюֈ����yt��Zo�����o�6Ѯ\A���	D�@ӝ.�����*��yq��J�H r��F�̮,�2^�2���&�����U5�� ��~�Ԉ�":���i�@����lS�k�W_@L}���$��Al�&C>a�V`b"1����I%(U?��t��-�ccrA�jʄJ����Lۂ��[I#� ��8v������r�L1�tE�4�ɢ�*�cE�#2iԕ�	&�ydĠ*lf�Gt.�JZ5�*gd�����3[�x�*n����� �vA��aH��,��oÌ'��ve$7�C�g�h�q\�#Q�8�y1[60�0���7�9����YT����:/9tn��4��V�!V2�A|�	�"`�Gߴa\����/qز��a*���Ij.b�c�� �]��˖Hɐ�a�̪�,-�,͛m$�&�\Gј��n�Jf���fr�p�TG"�ˮp~%@Fdv��Ob9�#1��H�&H�@��	���H�
 �ro@