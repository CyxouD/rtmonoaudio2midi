BZh91AY&SY��<7 �߀Px����߰����`<}M��©3�B�A �p�4M55MC��!���D  �i�FA�x�@=@ �@  S�h� @h 4�  H�F�OI� db � �����&L�20�&�db``$F��L)�mѦ�46�J����ؑI$��i|Ǽ��� �~Y*fld P���eD�$��`���xXCH���޸�g� 9Iqᰓ>P@M�q��%��AR �<ۙ��͐mѶN�;�Fb���q��]t�;O1)\��e=1En�$ �]�B/��¿G��lL ��~;�Wm��5b<����*oP@����j5Qу`�"�5�����ҍЖ%��pe�J�bb�L`�"(H�va95u"-%�F鋡x"��.Pf���-E�E#
�Q�����qP�xTe�t�����	ؐ�
w4��L�J㦖l�L�L��C����+��Zu���p@���h[ՠ�(ÇQ�
n�v10�N�vd�58�����٘D�D(\-o$X�(H��7j%��T��2�����-cux�q����+P6N$8�X�B$�L���VSk'�P5�U�U��b;q'B�q����5<��"���h̦�l2��6��LD��0� ��5��Ӳ��L��h�Y��R�`�euu1� ��ev���2���1u��KpؔԌ�)r�悍�"oD���M+�����Djf#Ra�����C�ip�-i<@/F�UZJ�;���Ec�sKI�"�;��ϯ����H$�	$� M�}�;���q�eV���Y�k$���`���a3-�q0
a��4�sB�Q@ �,,0����V��acUw�3cHm$�/�=6S�YK�q�L��ӕ�ڊ[-��&��R�B��f�N1���8�~�� |1ߏ�����Ԁ�\H�ٕ�+*����THu^_%��j?�=�-�@в݇xwѵ�ܒ�E���� 27��O��wZљ%W�W)��
]�:#Ċ�����f���M�� ,�&�'�B<�*Hu������nS�R2<<����)IJՅ�{)��Z%:��n����|�b�Х�ZK1�AGt	�[j�'�
��r9���**� ��y�3ZS�ֶy�k̵rZ%7�h_L+�� -�[��>P���Ҙ4 ���A�J�o�R�WF��}�'�`I-7��iѴ����tzʍ�1z��t�`��^Uf6  U~�61�'�>�A�TD���U�z����T�$�f� ;��8�_*�{�"ap��!��Ț,�TK!�4e$k);�����xV��D�24R�=Ѝ�$jj�N,��)�2M�I����@
������Ѝ  m ���6�0��w�>ޯ���}�/lhRA{yD>��okG�5D�)ϩ*I� �w#ʙ'��3�� ]}��g�gN7�|�8Wz�K �O ld��:��N���x���l��w]�8�
;�mcA���շY�D	$n���P X �)��]�4�̒�1��l��he�۞�,��P$�+�{2�\<���{�p�~;J�TVB5�6��� h�=��Q&0�Z$a�g�/��"�(HRN��