BZh91AY&SY�C�� >_�Px����߰����`�/>�� {�/j�!XI �=4�{CT�F�4� i�CA�~@�  h`�4 i�1 挘� ���F	� �z�h46��4  #a�5=S�4��f�6�M� �G�����ɢG���zji���@4 ���A�{"�d�B�h��Ze;_uT��y�@�2�F�3�+�Z�F�Y	�"��[�㽓N��b��v��w8pbЎ�9�t'p�ԜE��ZV��'x$�$��C��b�����ڗu ����=@l(�iP�Z���G[��H�t�Y�g�c�!V�M4Ԋ���������U$}s]�C������M�X��{��0�V�C�"�8L���e(@�&�Iv���|�l�ПS�a���Ʊ� �#D�nK�O�B	C��Xb�(b���w�����sc-B ���1,��&�.p�؄�d''l���4�ScD5S�*�e�ʦ��l�>ch[TC���*[Rʘ"f���.���q���t��a8��ma*Q�A|��o�Bإ�I4�I��`���Ӽl8E�4+`��8)���!t��]�3�9"ʦ�s�Xl?�ʒȫ1��T�Js����5�8n:��$5��eiz��9�f�C,����ż�H�C!Q"��du�y�Ob5☼�����/�~5]_9qF?<��� :@ HI$ΝE7��83z�wUZ���E̖rDV�:�fhƆ4r0P4,�`���L2,JG�b�$��3
��s:;e;/j��71�+b�,k�.�N]D�U\�2ہ�^iu�*�	��f,��x�z~ߏ�}R-+�U��o��4�G�ݏ�v��[p ����5������$Eq1��à߬�^d� ��m_��$a���6��IS-$G/�5���#��fȊ�Zs��r���$x��nՂ�!��o2�hu��6���J4�0ԥ큩q�ʒ =�i�u��t�N	��)=��'��ᐜ�|ҭB���Ϊ@�CD0!.�L��A�Z�&4��P\�#��rg*VJI!�%��&h�[y�yPd1�aӪ%7�����A~|I$��x7�݂��ބE��0L��g�)�FhTh��r�OK=d�se�)2� �������6� >ŒZ.���$��a�a�{l?����9��c����ծ
L�p��$���D#S㱽�s�`=���i$V��:[c.�2(����!@�O����H� �)N�P�*�b+��UM���&B	�D�S�� �P����|���5$�5$�0�$�ͷ)h����?Ӭ=S7�:���9ͪ��`�d�Ñ�bp�)=�I$6��1L=��,w����I\%�(H��'���aJ�*�����N���: �a��k�H�l띇�
S�"��|cb�n���$<���F�$�{I$W���F�e0��T�C�rѣ�h���:sI���E��U�H��у�r�]����I�d����=��[2�\HoR�`�S��w�]��BB�J�