BZh91AY&SY�g� �_�Px����߰����P�96�����:`�D LDƍ�L�&L���S�E@��    �5O$6Q��i7� m@� sFLL LFi�#ɀF	&@I��<PcJz�Sړ  ��Svڀ�H�	$9	�@px��������R�0la	5>������V6�,!�U��t�[<|��!.�<|x�E\#�n��嫣��]��G"p�U	��a��J5UN����A)�M�#;4�68�8Xa�l�ȟ��:[W^P�V�2B�d���>�/LBM�޾�[oQ��`�S��#C��V�k��!���3�x��B�/��**�ڕ��m�>Xƅ���-���dk�@�&:5�/:ݔ�!P(!�z��;�	�l�e�U惍�X�K������=Ir�3+����E���^�Q	�*2����%�b�&��d�n&�3��P^����vV{�Vd�#�\U�jh�H[V�^%3inUq��3j)QiB۰vP��� �5�Z1�k:�%�4��dd;�2����ѵ��̉=�]W����y�ĐH$�)$�	a�}=�<����c���n�D3nֺ����2r�AIAf���O� ��إ��TBL]l.3����HY0�a{Wx���b2y37�����/�i���{9ζ�Ku�O[݀��׃������4e���<匣L�Ԃ�w���5��bi��,]���ź���Y&�5�<$)f1�%}Y���荼C��̉;!�B[� fr��&��o<��H�)zӞ?��a�D{�J�۝|c��I�!(�R�1��P�E܎H� 0���"B���}Z�{�tQ}�XęZ6��:�zԲ,��ǂ��{i��&#�(�8 ӥ�I� �4v(�0:s.W5"s�]܉��-�j^4eq�ډL�M*�@��%){6D\�z�|)���P�!�R�s�r���P}[Jx/	KnE�ٔ��|h%LY�De���E��W!��J�a�a�{f>0s�9���i9ػ5	��MT���n]�����M���@�|܋�l%��qM�Lh����v'��������N��G5�
�E��f%�r��0�$̀{|x �����	b�}dh6h��(4A>�C��I�t���_OA9[����fE}�0Ga�ٙ(���ߏ8#�2_�E��5��Jz�5<ߒ������v+ZY�z���r��)pE�O�nK�5�[cbk��,h#�،ukzT�T��G����J��K�q�r52؃AЪի+�{p��"���Q"��v�&.	�>������Si*5#����\�$%C2;�*ؓ��of59��2FZm�&���"�(Ha3�}�