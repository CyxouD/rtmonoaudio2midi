BZh91AY&SY�Y�8 �߀Px����߰����P}ޗ{��V�+N�$�ɢi��xS�S�6�C��OHzF�='�Ѡ��)��h��4   h S"#SI�46� h OP��M�h ��    �@@@���ѓ*~����@0�2!(�� ���0	��(� ���x�d� ����q�E6�D"�(��фEX�.W�{� 9Eoߑ(�1���a[}b��YLjgv������ٺ(j�T���s�'�M(�Dl�zО����ǁ����iZtA�Q�� 'lD�H[�˞�Ӟ�� ��7�����u�X(�6"M�2�r�V���X��sE� ב�<���$j�@%	E�.b�cM��,���Ŝ�oc[K���A�҉�p5M�v��؜+���i�SEU�c����o5H���,�-w�QJʂI��Wu��X���޲ @����r�f�Wb��[Z���J@@���Eu3b3�K���pzN�HHIz�I$
 ɾ�^'���W��ѕZv�tJ8۵�nQ�'��\j(��5"Q	E(�/ ��f<�q���S�E��hI��w������yJ[=W��pZ�vxJ����W���㋿���P+)�J�Θh���y��r%]��H}�&.w\'�ч�8�Ξ�����5�>�.����]{Cl[�?��-����y��r~޾�:&�$���_Q��ȮF�3���8�6�� W�K�͸F-B��D�
+��F��/V�n�%���=�*����z[4�d�7(u�}�38Qb�2> $+[iL�\�GӖ��D@�lΙ�ҽ�e���߮�E7���֪)/�@�z;�v�vG��u�]�& F*R!�J�n�J�u�ݬ�����X����Z�%��&m�5������\�S1� 'f�61��>��~3!|���<Y�z� ���H� yp8�/ 4A3��������R�(����cE"C9$�FƄ�	�����V(� g��M"�g'h����A�xr��(� Ł���	�r�Ѝ @�ePw��f���ه���e!�&}�=%�sc�Va�5+Y# �o4�=��� ���qL��D\x�~�
���ȯ����rЕ��b�8Q��!�VD�P���"��i�$����ZD�aK��Q�f�H�7a�ʠ� ��d2�M��1�,ٯ�Ю�d�{Ya��I�{,�T��&-���L��W��j*�#�\�3 ���1)��|m��cS����$f�v�_�w$S�		՘��