1.594920634	New Point
1.995464852	New Point
2.400362811	New Point
2.813242630	New Point
3.196371882	New Point
3.591111111	New Point
3.989478458	New Point
4.391473922	New Point
4.838004535	New Point
5.181224489	New Point
5.381632653	New Point
5.579319727	New Point
5.958820861	New Point
6.175782312	New Point
6.386734693	New Point
6.754149659	New Point
6.781587301	New Point
6.968888888	New Point
7.196938775	New Point
7.553061224	New Point
7.585714285	New Point
7.612244897	New Point
7.782811791	New Point
7.996734693	New Point
8.363990929	New Point
8.401269841	New Point
8.569523809	New Point
8.775056689	New Point
9.150113378	New Point
9.176961451	New Point
9.376507936	New Point
9.578571428	New Point
9.975873015	New Point
9.999092970	New Point
10.200000000	New Point
10.422448979	New Point
10.765306122	New Point
10.787482993	New Point
10.979047619	New Point
11.200000000	New Point
11.572970521	New Point
11.778321995	New Point
11.988775510	New Point
12.348662131	New Point
12.372244897	New Point
12.583764172	New Point
12.795646258	New Point
13.169387755	New Point
13.200000000	New Point
13.387755102	New Point
13.598185941	New Point
13.964761904	New Point
13.986031746	New Point
14.008163265	New Point
14.178684807	New Point
14.394195011	New Point
14.754965986	New Point
14.775918367	New Point
14.795873015	New Point
14.977551020	New Point
15.184489795	New Point
15.566122448	New Point
15.585079365	New Point
15.787120181	New Point
15.998548752	New Point
16.343356009	New Point
16.365804988	New Point
16.384263038	New Point
16.571337868	New Point
16.764807256	New Point
17.133560090	New Point
17.158503401	New Point
17.181451247	New Point
17.354557823	New Point
