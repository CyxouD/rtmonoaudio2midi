BZh91AY&SYz��l �_�px���������`�M� W}T�U�"�h�Q�4�2Dy2h���L�J hd  �  �風`�����F��F�2L4��%4` L     F"Q�����4�F#a�&��M	4�hQ�
zi7�=M�0��a=G��
f~<�)�
TE!T�c�~O���?��`� �A!��fG�T�@%��M�
^z�^O�J	e.;[!�"@A���S3�-�6ғ���`� �����0�p�;)ݒ�Pa�(,`*�A�Q�$�s'Q�R"'�%�)(A��eu���^�CR^1��_* ������ϏV,($DAxn�����?���'7��:&�Km/qٺD��DfD�鄶b��!55>Bv��([��TY��첗,bH"��M
�_cd?�R���Lv�D���)�^[F�nSd�r��X2��N����)7q B�U@]{�)rQ�R��;����0I�uWD�g�i����[YsI��*��c�;DS�(��N-��1a�Y�[~S�lX�ّ��Z���f�PF�B���$��]\�d�K0�9`9w�ЕR\�(Y�"�RI�d;D&�k������P,ݥ�`�Ն�|�-�$P�g����qͥJ�̠�̠"mDSV&���2��'K�wV���Sg�烉i �� BP$�R��Zz�/��쳅mN���H<�6����T!V*$�hJMē��
� ����	�f�	��=X�T�`0T�z��hĀ��˞�=uOĪvY�ӣ6�!3y�p�HӘ�/��?U���'���g2� 6h)aB G�m��̳6 �2���S��Q����A�ilWn�{�y/΢��`B1Z5���}H.�T�H��n������z�2$�^J�Ȗ0\Nɣ�!*o��j��i�@}��g� E~iI���p�Ӛ�[�h�fz�-�
Kŋ��=��q�=WNq�j�K��9<c�7O	`��@i����+2O@b�ʆ��]�\7M�N����CQH�qNY�3�O��cރ0�O?e��G�����~~�ȶ���fH�[����@"R��QG��)�~&�[B�y�ߋEٙ�.�Lu����Pj{���#r�=8Q��HE�����g��k��ʽl�t�a �Ɉ� Gw�#K���8���L�Cg���f�<�0BaBu�b�2�����5��Ac�HA�粙-\"l�4d����4��=��D��;�p6��<� �T���?'	�k���X<{�q�;�7w��� ��߰l:�-#��<��ԧ4�G&��N�
D�O@pr($��^�;���Xsr�ŝ+C��,���%�ZJ�����.x�~4�P�������V6fwj��~qF	>��E�PKi)��N�����Q.��mU�k��B���Ҁm$�M����巠���^�l�QM�f�\Q�?<� B/G��Q6U��-�P�F��Fˡǋ4�_aw$S�	�f�