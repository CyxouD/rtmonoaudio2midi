BZh91AY&SY$�� Y߀Px����߰����`��M� �8��@��I!O(��F��=H2=L�(2O 
U=@ �4�� P�� 9�14L�2da0M4����%2D� h�2h     9�14L�2da0M4����$H��(�����='���M����	 M�R��! r�P��$��z�����~Te�T@&��O�'s K�*����EX\��ηqՆd�
ˤ�ٌ(�{=W1Yf*�jb�5f���bP&�"���Xjk���\���?���f�%��Z�!�W8c��¾�$1�dbF�S��1urBRzH�xtW��y��0�L���}�������nf�bV�����Q.�'�D�wS�n�kW"�1Wk��Ɉ9�z߀��;`���u]D�l�"wAƒ�����Yyλ��G��������ռ�4^q�>����t�K2�-��NR�fR�4M���&+��cɸ7S��钔���Sу���7 3]��9r�]��C�n
H��D�/D;�݁.�3�q�PZm�4[5[;48/�-����m˳ʢ�O��K�% ��L#2�G2�[�5A�];�Y�Y�0��R*F�/6#5�6(~5�0�ӎ�-��db%ve��Kg��go�}A�R��r�lf�;��p�t�Z+S����`����}�@�$�AK}$�@� �2l���LG7
ŪVp7b%�ֱ����b�p�1��ܴ0��� b&���"L6��Qa ���P��7l�^�Ʌ�S�k{����X�������#5tf���e1��z�G�)���zC?=�e7���Os�{J���D@+����Qe��1E��.�I9��z�4���cG��~���Hr��M|C�ͯ�?�K؋á�� �@�/_��G#i�\"	Gb��!��_9�x��k8oԿ���<�� �Ի�¡�V�ңC�$�'�_�t$@{\�/�k���J���֔���3�cU��s�P��ZڮZ:��A�D^@#��N��F3�}0T0G��B�"B9bWթ3K�w-�H4�c�I7�������� ����P�k�f�a�� ����Ρ:5�z��sf!�?��}DಿՉH���y7��V���j��]49� ���61��?͠�(D���L.�f�V����L����_PB6���s���`>�tE�h5E��KP�+"3&�I\�HP/Y�%Ou������p��7�#\���(�PD�	UD���x�B�GgO��O��3j9�@-t �]ł��S� y��Ɛ�ű�� �����n
摴�q:��b�lb>lzP���8WHk� *vVU>�%�����˾��id/ZSX62�A�fN�����<.�}Q`��} ���9H�$�Jed��8Dy)���[{
�g:�I&2Jv �s%VYLgsOC^:1 ��A"Z���=K_~���1���(�܋�4hpm�@*ّ��I3��������&HƧehQ�rE8P�$��