BZh91AY&SY�,h� 	�߀Px����߰����`��xx=  '�U�EI	�=	���5Ȍ��zi='��MSA�~F�R� �  h h ��hhhb4d @� )���h 0`���	���dɓ#	�i�F& ��#U?D�H~�S���y&j � 4���"����U)eAB�(�PF��q���A���f��	<@A� `W�A��
#�0����K��=\\�\7�5f*�G�5՚W�f+)��J����'TP������r3	�(V\�Ka�FB�N/��!`�,y�����n%�T@0�uWA��:0��ǚi�@�����і]�� '���;Pv�,��إ���e��h�NF�%��T�F	H���J�q]!e@�ڄ�BL�
�q:��9Bd�ې8
*�� �늜
��q{�{�4nk���*�mdUdA�{v�p����c��t�¼B���.��jN㙠�j�`�^�@|-x1U�8��=�!B�F��c�KH�����(�v�#ME�@��"������M�Ֆ�M��UYr�J�Q�ʕ���LV�ڃ$�8ڔ_C�a���]@�	E������ �,�X�Ⱑx�4��D]�B��
�+�/I�0�$��y8�O��3����<gm�EAr�flN��|J�N��wnV�d<�V¢8�E�lEt��mL�\���	m��&F��-�nwzd�XH�`ӷ|��}��Xb�Z(R������rm��P��m�o>�췑Q�*f�Rċ��θ���D!<_���i�Ȋ-zG�˙�s�����QwBb���C3:�����ڜ��H9[\�T��Dc��C���ؠ�[�@�u�^tU�{���*�ʨ��W�Oi�%��ˊ�`�#�U���=z�a����+Yt�ll�Jgb�^��]�0 S��"[��X�"�V��(�]u����#5��Tͩ6�S��#�p���.����9��)������}�1�!!%��I P�Mx�"z	�ş�H��OẢQ��*T�%l�

��P�P-$�+C��ЀB.2�`P��@A��wm�P�u b@�7�;�4dH�6�����e�y�v껉���wzuBy~�)����x�>�(��k��.)½� }{�W���3�z0���0��_��Ǿ�F������s�M�V\�d�ص�w`vI�a�9u�A�@|i Q��������[�_ܺOd���Ó�y�m܀�O�
^�fc�k'Gܘ7A"8����u$�-�_���%8'q�R{�VOލ3i?\!S'!����
���kȂ�(t�-B2�ʦ��o5_4�l?����-@A��ÛV�1�M^N�5$1Ӻ��'�fa�L�[��h9�{C<���uXo�02	�Ng�)�Fq�G�!P�8u֞�Ն�ƃa-~�pŭ�9��}�L�/��
�ka�a�{fy�먥vzx�<���F:��|qQ�O[��O$��8J�,���H�&�ÖX8�F2�MK3��Dh1�V:��B�Q0�#���H���ȵ:E�K� ɬ9G,���h�)�sې3�����8��H=yj.3�9j.�9�=�=_kOAFk�I����HO,S�Q>É�и��ϥ�a��p��l@@����$v���m��ա^��Z��У�� ��g��*: ��Hi�Y�`�3��U�8��%��43�ֈ9@o��Z����q(n%�u�u��k�܃�1�$��#`ܗ��^p�~��3�"6�)�t�d�����fG��U&'�}5�c����&H��uj
��H�
E��