BZh91AY&SY�nL� �߀Px����߰����P��M�9�@�H��Lf��!4�!�H�����i�jz J�   @   I���$4dd�h=@  �9�&& &#4���d�#�2��Ěx���z��i�z��0�O�ؒJ�H�HH��H�!(�=�	?��R�
�2���'��@`0E�>��(��w�\<s� �ٳ�Y??kX8�qX꺲����]�.�V5svͭnG ����F3��G�q����˒Zc��A!�dbG#T�7��G��U�� Z��;i��z�`$�cOw��k���\�����2���[�k�H��Kr1��T��D������Q֛#e�87���ұ���@X��H���/l�ܙ�h܍�:(iU�\�5ʩ�gkM;��bI�BѨ]1�2�7��.�MmhR	��TE���@,�\R�QtT�Z#jj��J2D��6�0GȚp=�3�[�p�����"h@6�j�Y6���0��D�2EP�61gp#,�%�5$�k��̗�ڂ�ʾa�ǀec�J����-���~�|ÒJ(��UP`IE�o����������,�ʬ`�3yj���Pެ�XFg{/`]��P�1��	1rac9N
�L,���\ ��h���>�W�Z�M�f�yO����S�v�&���)z���L����D	���H[�����MMha��u�f��G�f��ǔp|((z�{Nӧ�!S1r�-2O�e�������KԄ�����;��ܺsE�_�Q"Z\��tA��®Ku����>@%�b�ƙ�QD{d�v�I?v�f`�(]6^}#��J�Q��R�cn�.��W�%sPӌ���p4��d��4�;$Ґ4�u�0��tSB;L싋�D�I��3L��L׊�2�y�&�0)��kא	^]��n�F�|fDV��&R���H6)��S_PL|u�`�Z��E䥜CD�n#/���":�W'X��Eݳ�so�[Oo��S�\�Pho�@:�K����}�^�(D��r*CA�$Vjd�cE$FDӡ+4  MKι0qe$���ܑx�����*�j�A*(�9�W�P@�+�6�T��J9�J�Ü�^:
E1g�y�͉gқ2w�Nx���^Ѱ�]-#Q�8;����JE��ð�2N����(W{�*_�1�����Z}�as0 ���I�0o#��k�w[m�h�'�5[m�W�	]v*�|��`�"��rz�W��9�=x+���R�C�E�͢׆�w��k
���E1� |�+i3�*�d���q��#�eE�8>� Jvdo,Q��8h���3��k&H�q�k	���H�
�ɞ�