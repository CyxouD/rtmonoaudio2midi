BZh91AY&SYkɂ$ �_�Px����߰����P�����W8�:t	$�2����F�h�ɑ� 0A�~�BR� h�  �  	L�54�F����0��@   JO�4i�����6���  � "�	���S�Q������`�O(�R*B	h�HX�O��|2��I��H �4�K٩B�H�y ��!3��)Ha��{=�ҫ���꒏�R��m�V�R�c6rR��I-�bBvm�8��I�26�m*SI�&�X�֒'t���Di�y�?�q�[$F\ĝ!ul�3CJW� )|�G�;t��q�1�����=�a�ȿ��{��}Nof�F�2�v[��)C�)���7��p�}̃v݄c�e��.�#���J,#�P]D���u6��-�&�,�gwSN�X��P�R.��^j��6��v�r� ��@F�my�V=K�qjhD;�ș�  H �S0� ����S�ք�ةX����d�)'r��E萶 ���V5V�J�	2e�0�,pS�[I.�H0D\�)�-��O��f��0�8��t_L_Gh�-�Z��� Î��{�MP�%�>��?�7�����$�@���6pD����-�N��D���X�.���2�%�	߁*���8D�R�U��i��⦅�U�A0E�>�l`�3!%m�.i�w4a�FY�ϒZN����k#����߭���xl���oֹ�>E����-���M YaA|���t
���i(���Zl�6Ϸ,Kٌ 2�ۦ]������FZW�� -Pnv!�oZ��p��S'�r�8���*a-�5/1�@yG�K<v%��'%u��Z�F�"W�v*�(�ҙ�}�X�r&w��1����۝;֕R��_[�[��e1CD�"Q"� l|`H(V��2�W0mpn.>���I��=:��1��y���h�W)���_sF���U����]ɒ�L��`  '6Aa0ɪ��Mm5��7CB9�)���D&}�%�c=f�)4�^ƀͥ�.[P�:�`$��9Xfi�؞y���E|��l�3ڤ����U��7s���$���;Q9%A���Z�@ohT�'AB��q@�!�~�1&%@A[k6$t�y�R��N�w0�@���b�x�  q`|>m���"I-	$�q�AɆBB~�۽Hzs�F�良��U-f���O��8VH�9���&�ɦ <�[CQpF*��I�  Q]1��x����\���M+���*f�����} �4��&�1�,����#�"���5Ur���KB���i��Un�V�I��W8�0I����yR���a	���m���c�*�m�\��2�k��rye�BJ*�#D���ǀ�2;�
�1���3rF�&H��r�,���"�(H5�� 