BZh91AY&SYjٱ F߀Px����߰����`N�-�9�1BGfR�
m#6�4��'��!����bS��bi)  4     ����OD��F��F���b4���	L�T�����4�i���h�� 3P9�14L�2da0M4����$H�4������mC)�l�A�4S�� ��$�	INHH�@�7�;�tF� :���#,����Sdx�HFQ����4�0����p�Ն` �1m8%�0�^�mb��VS+��Ԧ�J<���
"�J�����$�*+T�$���;
����c>t'֜e�$Fl�e��u�{Pdw�$ +KHHKxbb���rL``���E�vٰ<F�I�P/	��>�����h��M �C�{g��@Q�w�
eڜD:��}""˱��� N���$���'��Z��Bݗbu�n�5�v�u��lcp�V���g1uo#.��
�:mr,�·Ҍ=��1|a��B0έ��䝤`c'1X@�1�⠢�x�M�;`ˌ�'8�Bh[���o8XU��I�_!@LZ�l�W�A�@wX[3�as� ыhz%Ĺ���P��p���j�*�\�|�E�A��:U�}�v�R��CR�e1�x�,�+�.c���K���fjآn����{�	!!%ʒI Pd�kn'��{�8m*�z�o�j�3��B֣)�`I����IM��@�0!��E@@���S(;���U0�����mi 6,ř=�@JW/�M�t�bΡK���?O�R�&�UD)�B�;�_�ÁFJ� b��<_,Dy����x��cz��ң��2*f3�Ab��~M�M���CC` �!p����:��ǚ٩%o�D�l��=TG���[�W�3w���
������s3j(��$i�u�+���1�(^k/���%('l�i��f*�+M_�r��1���8m��&
�BJ ��;�#�?Dv�`zr.W5 9bSv��,W�h�f1����M�0)��׏`,]��8�"9H��ӆ�K ����nS�8�j���1��Cl��qc$��$��AY�D�1Sq��>��n:�� �8�a�a�{j<sm���ղ4Ks����֒� ����T#c:�=O��"a��A܊�h>}d�}��ZƘ�Y�4�J�D	�}�А��ˋԓ�g��䌈؊�����c�d��B�z��&X��n�&��IZ,pj�S �� ��1�yuyKo����U3(����9����9T��!Σ���+���@�I�p.]!����IP��+�,fދ�Z��:�Y�
1� ��Z��# v���)ۨ�#>`�D�>SK��$��#%U���
�8[7�� �3��q��Dh�R�c�E���`׶�=�_y �KY�\*u�y��&�hX�3�a�-����E������.Q��}���c��OH�ɒ0�v����)�S�͈