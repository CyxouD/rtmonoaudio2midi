BZh91AY&SY���g �_�Px����߰����P^9l��7p�&t�$���
~�����)�=	��D4�ML&�E4���6�CA���z��0��! �ODh�d2z�@4   0&&�	�&L�&	�����~��<"x�M�#�  �����*ĉ��h�!(�=����8|j��6�j~$��u�!�V6���*�ֹ��g��B[d��I&}�uA�~���Ss4��n��+�v��f�c��LQo�F�����Պ���s��׮3����H2dS��ԃ(Q�� Q;����y�����2&BL�����6,\M��9^��h��vc��:7�R��We�.�Ɍ[Uqm�͙6y���f�˓2�g:�*s�n��c4lz��T�TLDDX<4aA!t�V.�k0u����:����*�J]�H4,Ȭʑ���.!�ɬŪ�,j��$��$�����B�	!�#(���D��]kq��.*�i�=��Z�rH$���$�
�w�W)Iyx8��k�bL2��K�E�J�Z��c#kD|5�P�͵��P�#�!����L4j=ʖ��&d��P��w�Hq$��m����g;��?�_�������,d�3\y���ȥB\�ק���Q��"!�̓�@{��������5�h�鑑'��Y��7��A��ԋC���%�!p�8��=��^���#J^����si��.��b�Õ�|	{Д�)u����:�+zDx���/��ݔٸiO���,��ƵU�c;�/EFj�Uv�;��3��iGd`&�TN0(t��/��ClW"9��|
E$��YJ��3�7��0����M�^V��T�_J��opl�F�~fDY]��$�%�H4�ڍ�Ы�PL{���$�|���3r8�5�yC�f8Y�!�+����D%��fj^՟� ���xi�i71��e�K�sEhK���
\���c[X�`�>0wFH�o��X�h�1D�,�
шDU���B,.h�8�Du���Z+,�uY�(JV�o<�	�IE:���j����HK6�6Yx�(��|�N$�8HY����')s�:���_d����xv%d�Г�(#�2N��A�BP�ପy�4��ϲ��R���B�d��5��N�9����<�I�'�����,.���iߐ,$Tח��%sBU˄�C��r*�B���̱c�[n�n��"�I�@r�H�Q��BϤ��+�fr����)���289D$�fG�R�IÝ�q3��l�"�c�nb�Q�rE8P����g