BZh91AY&SYu}} �_�Px����������P�� q�S6&Z��HF�@OL�����MmCMi�M�5=2IC@� @h�  ���LA�hb  �M40&&�	�&L�&	����)��b�OSM�OCjOI� �< (�p�%a"  �$�a 8�I�"�$%��r੘�li	59���HT0D�mL!�N�޹8[Vd������~`��u�n����J�8!TT��,��j�&�.$i�WSCr���~�s�FmQ#,�F8�p��	�A�C�j�k��A`C��I%<��b�5ϻ���Ji	6�y�uێ}a�O��i�Ղ�`ߣVwr�h>F��%�z�E/|�Z��1YGY�Q�� �Ai�D)���D�`�K�vu~��[<nٕ.�v��f��	s,�3�f(Q���9���%0�[fE�����"�CH6���
�M�LF��D3���%2։*�],��p�D�,���"T�Q�B�ܺJ]���	o,�Y\U�m.������ڳ�3Z�X&^!��,�
9L��w�B�P��Rb5�Ug6����[�Y���~�|ÖI�߱��`�%�[yO����ᵉXaW�1�%�QY]0�2d�q1@�����؉��		1q��H8�u�х	�-M��b�EmV���ꦏ9MU���5�%����w�?�/������aO]?p9�+�Fu:B\0i���(��	-�)���@��RN�_��JJ^���m�v�V�\	,�׸7L߀�9|8jd3HK����t	�s��:�Q2Y{TH��X�3��t%�^nU��Bq7ZBQ�%����N��"NA=s�U	�$˳9��SA;eQ��:�.������nMKP�Ϗ����P0!�in�)��-)��rlT� �R;�g��	�$���'�jf|�&u�a���n��oA-�T�Ԅ�$��7���:�ˣ*``I=���ȡ24K�K�Ѐ��m��JI�s⸜ˌh,]$���P�|԰G���	IN6�wI�� �e��5T��+Y�2�X�$���[����Z�w��# T=��E4�R2�d�6�4c$l����Aj~�"�e�)N�(Gj�3J�.-N3J�A)�I�N����)�0ƀOW5�Ƚ!+R��"��6"�CD)� z{��bz��9˽���X���xu�6E��i!�1�^v*r1�%w�N�F����ר0�fHI�Ni_)�Ȏj�7j�5Jԫ��ք�d�A_��0F@o������z�D�9�8���1CAs�'f��,@�=mlR�����s:�Ո��'�qX�%VYLӆg���a��$KPٰ��T�l c��C9��^F�2�ȷ	}��J��T�2��.96m�H�i�aa��ܑN$_E�@