BZh91AY&SY@2?	 C_�Px����߰����`G�{u���A ��$�i���=2���DSmMh�L���	�*    4   T�L�4h 4     �%P�hmC@ ��h�sbh0�2d��`�i���!�H��� )�Jzb�Қ40��! ���0���$䄈�p�n6�@yz�A=���` d���f��B1"�6��,�������s}�������أP�M���qR]%) ��h-�ȐP��bd2�!I���B�O���!�$��� PC��z,i��f,�̧��Jmk�Pf;ܤ -v$%��PC��ݦ)�@�w��m��
�FY<���ܼ: ��ڶװ�&fik��nTH}���a[��O�!��c!+Gm�� N��f7`����U�Pz�N︠P%�#��X[>���*.�l�|@��0�b�Q���V>��,5j�@t�	I���F�A&�}��b����45�rX	�t��A�⮙�$�j��b�;�+��\aU'
`�h� �8Lt'Xץ��R� �U��vXX�&-�8Z�P�ʣ�%����6Z�X�%�&ڞ"mC���Y���T�CDP�ِ�&�5��S��+8e������$	=ĒI �:y���#��tE��֕$�n���@�l%�$a����1b�U�dԌM�g1@4�XUg���T,Xa{U�63��$�Md�{=��n�3O?=�q�v-su~�e|n���g����j{�e��YO����.=zm���ʁ�HU��6��^?J�:�e+�Y�{�o56Q��=�ͯ�į1^Z��]��y�ΝˇDJ��*<~g*�N8��t�c�=��1g���[�/ќ������tJEy�+w��DQ�k����8��į����i�;��[���xf�j���{iA!�X`��ЦH�A�Z�&T��P\������*5V����Eܚ&i�oE��F�e��V%7�Ļʂ�|�A�_ ���/�Y~�@��N4��&$a����`�|T��Y�1�ϿyA�=�6�R�m`vm�9�v��]`˅��{%��?:�8o�\o�fܖ�s	!�����'�c��\�(��Qbd��T'[lcE�F���M�D�<%Wۆ�DPX�Jp�B6�#!^���*�Q�2M�%�Nˠ�����M?�k�*7���A���9��c�}e^�X�"j�veK�RV�5��f��#��z��ZX�@���B;S%��i�ր�ˊ�>c�aj���ΫJ��~@fzN~j��PsTu�\��Š�7F��Ek��XZߚ�Ҹs��\t���+�|��>LUe0ђ�bC�r�L��6ra����80�
F�Z^ʕ�P�3����/��)�\�2\��=
Y��X�����FcS��k&H���	���H�
G� 