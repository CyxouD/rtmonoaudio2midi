BZh91AY&SY�Bo� �߀Px����߰����P�8� ᎌ�cj$�L�Bm4�%����&#)�b4�jSƀ�  d� M   $Bje2d=OB4��h0`��`ѐ��&��%b����S�y52P� p�� �KT�(^t�����~�B�~�X��ᐳ��@����D�H��/��n;�8eAvU����~ ��]����+�ٔ�����2�*aI��Zl������?����v�*�IC7�V�8�p�h�FfͣITg��X�DC$�TlɽUA�w`6����w�� ye��z�N������f��v0c�����s���8J�$�
yF9x�QL��)���,�p�h
�ba6���u�O�}D$}�veȬ�$9CJ��o0�Yqud�{b*1��h`sX��JɂN��8��*TZ��g� d����:y��Z��J3(�O����ꔓŪ�#���h����l�21Y2��lYK��	�$HuB�%QDh���YAB���{����^�i��\�e.�\qr�9h������66��ߥ��`�%��1)z:Z�V�qd��#+�@�KH$k���H�͟��T���84�R�^Z`�1�l00ɫx�oaf[*������˴����7{����~�Oo�_����q��~Tu�ӡ���nS@��ٿ���]�BLU!���Ƃ<��5��eWq��H���"��n˴6�>a�(�����"���39q���9������P�����#�����te�ט�����(��_���N���D�ǲڀ��r�5���w_�JpN�R{�'����X�٫5w��l��h����]f��5�JA�ke&�A\\�F�A��Xj�)@�>��.L]I.r姨E�1*���kʊ*�Z��s ��N@ՠtע�6��kV��Fz؟4gF
�1��C�4���L>�\�F�Zz�����ߺ�W��� J5�a�a�=�<����zxF��1vV+����� 6�G�3����(3 ;#4������Ƌ��N��Ā�5>�j$E �)N��F�4%I�"�%9&Q�R��\�A�@��k�����̂��A�-%P�8������6M&��jV���9��u����D�f����-K�h�	������ؠI˚�2���"x�Y�fq�hJ��5��b	8vZ�!vQ5��d4F�ɰY�v��R�q%c�ؤ��;i	�(2�֡Sd	F�0.l*QE�9>C�F�B���Hh�`��xI'�	X6�	z+~��hڙ�2�iE�JnF�v�?XJ�dx(ɉ�4���(�x�4�'���ܑN$:Л� 