BZh91AY&SYA��� �߀Px����߰����`|�-� ���h&HFA5=5Oh���'���h�OSCj&FM�5O�	�J�a6���0&a1`LM&L�LM2100	�'��i�z��i�@  � 9�14L�2da0M4����$P	�dh�����d�F&�JB�.�����i$�� ��$A'�=��ߎJ١�`�p5d�\��BI�F6��iaf����Z����g`�~a��u��;KT;���x!N�U��-�P���P�WvKd*���9���͛N����(f�Z�1�wy�#0Љb*�,s��܃ ��qHV�DI%X�Ts���I& C00yh�:�W.���n�M�@�7��I�*�uu�"�f��`���s�FX���fCQ�5zzGVEoĐ	�ck��$|B�p	�'\��lg$NcN�˾�в]C�\8
�j�G(�i��N-j�;^�O@t���D��9J	���`*�
����b��`nL��q��t�Á2�1%�;�l<;j�PQO�N�UAñ��bɝJf"g�FP:Z�6�cL-4s�1i��uHbU;_�أ���mݴ��a���L�����1bY�9��f�i&ɗ�w��e.V�7�k[c/��8 1u95�6*4Ҹ��6b��|�~���66�����D!Yy;j�JK��Ņ��^	2e3�L`2m�=�qF�ؒ�$�%m|���Cij� 4�Uc���(,XTaf��[��T�LV����Q��4���f��sGoo8K�t
��7�ƌݝۧ,9j�Qk�XU�F
@���综��P���"et�{hO����2#�[o��χm��$�Gӛ�k�r+�Vv����`7��&���iWX�%.�;�B�'�9b�!�G\��1~9m D~�w1�Èi�:(��f֮�T��+侙�ٰJPN�\b�Ы��-\h��A�\7��K��5MH�!7��i�4ѝ����<f���~51Pl�l�3;����$�ep�NM�/)}ʊB���q? ��(|"C��7kL��o"�Ԭ�ާ���0��C�I�d��.l�`R\B�c�=aѶDqZ��I�q��,lc�/q������;����,���C9����3�8��S��q�$���R��i��Ѷ1��!�$�F愑w�S�]���'���H��kC�Z%(KVJE��W�A �)�:<*	���p�����"�^�(U�0z|}%PtH����T�k�ٴ��6k���dQy�ϛ�� �ɇ�ޙt��@|����������cy�^�޵%�uYe=@�ɥx1%0����ט㖓���0�'�A[m��0#jSU�-,/(m�'@Y�"x�a�,�fȩT���Qg��-��[(�HxE'�	�6[RޫZ8�Bն�r�����J�#-�8:��F!���h�.ݽtٿ"F��F�Ŵ��ܑN$f���