BZh91AY&SY��]� {_�Px����߰����P��x��64fe@I!'�M1���4�Cb2jLhJ d4 `M4� Jd�&������4�@�   ڪd � ��h   H�@�i&�jQ�i�zM  �"A] @�����	( �P1�m_�B���4ReLL���q(@]��Q����EV׃�k����(��pJ?aen��}եCT�Y�m���⵶��\cjU;%j�V���9o��'�Z�;��(�".l؄����#s�1��ˍuU��)V���� ��9���v�֘!69��Y�j��k�u�^�d�S��:�:JU(WY	L��K���n3|K�z�SZ�P	@��p�� �Z](�T�� f�|6g7H�88���3��UT>�(3Uv�R]��	J4�D�)E��Pمc��1&e0�� m�zj�,��YM�RCe�XG̳��;^^T�&d1�R���E��
�5T�9nlXZH��P/4�6�Ց��iT�I�Mb�Ԍ�NZ��1j�uB��g2�����|�y�66����(#M<j=��^~��X-AV��(��3� �FQI&� �c4D��@�L�2TDko"9Q��.N��aRa[S�43 m.e���{!�(�%(��mzu�o�'���e?]ϖo��_�+?5xSc�9x(�)v-?�OB��k�i!]#߀�f��ه�5%/Zh�q�7��l�t!dWwjŴ6ɼ�q�E����B��@�w�O1����KN�Vu�<~G,���9�M\7�a��Iu�|�b������#;�&�'���B��=��e��um��*�^��R�a�&�.|��oX��;�����c� �Z��U�nP9ڍ��11�6�N7Ղf{
�י�Kz��)�J[b���o+	����!�U5�L� ��q)V�tҩ�PH}$��K$�q�y9��:bߑ��cd9�?
�9m���vlc��xA��ղv׽��̙�C�l�b� ���.���b��</���\=�抈4xI"����cEQ!�$��� 
'׍��X\�&{\�2F�h�w����5Q��� ���Dg⨱�`B��E&��b��S�0n��*C�#WK�OAK5�soY��3
��1�GI�ݖv*��O��mL���s� >0B��E#C�����M���jЕ��_�Q��!�R�՟=�ii�7ʣ�
2�0�NR:X)�T��S�`TH����*�
�T����gEl9>#�#@����Ne���:R���F
��`
����t,]T3�h�^r5�)܌��;`�,#2;��h�/;�{1��$^ɒ4T;����.�p�!
��