BZh91AY&SY�!` �_�px����߰����P}ޗc�v��P%�����!=	��(�lI�P 4چ�SL�B���m@@  4 )���� �C��P�i�#!��i����        $M&�����b��)��@I��4���4 �A!�!2���a� ���^) H � 4?���DB0"�m!�U��vq^��^��*���d,��:�qcx{�Ly�>R�ͪniK�9C��T�;v:3$������|�B})��Hf9�'�1�f]O��G$�U��AP�i���v�& ���~�sf�xu���Ť��h��nhNN��M˨��x+^�2`���(�Ķ/�Y�Z(J2-�$�V�q�ڬjseb)�� ���,#�٪	�2�E �DTp�G0�"� �h����ҤM5����F�Y�)
��H�N�N��fQfT����I1��JĂRT�X[+'7.��ru{xM)!!%ƒI P �M���x	��ǪхZw[�%���A�W}H�P� l�r��(5(��p�M� Q�,���8-�L,0��y��@b�fOOH�e���̛�wxanLYH��-���~�㋪b���n�l�Mf]xqW n|��Mf�~������N���� 4���^*xUkw-@.m��������+&����]��<��ñsf��.�<"F�^3e�<g�G>u�˙�\ 
8���j%l�t]����7���:�%�����	J)�UE��T���&��BfN���L{"�#sD�&��=RiHs��0�A!Ӕ�(�H������ �ߢf���5����e��I7������� �����Q�S��j`���T��&�*^�םW�f���O����$������L\1[d��B������n 
c���=$����hD���x3�*y�/9�I�ڻ����`v�.P�����z�T%��-"3&�I^Бj_M�$"`2��I�3�p�E�MY��J�A*��9���Q B�G{�y#`� ��Yn��b���@�|��bW��ٱ;���:`�V2F1Ѽ�nΕa���F��ŦU���h ꍒ�������o��Lı����c&��n$�0o#�����l�
浇BC���PX�U���`p&2*t߭� ���Kz{�Zћ!J��2��[z��yH�P��I���Ix*��$K#�p��Mw֨Rte�]s��
�d{���eߖ��l�H��H�wh��H�
 �d, 