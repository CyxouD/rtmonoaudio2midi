BZh91AY&SY2�0; b߀Px����߰����`�� !�ATH*H@Д��&�К(�F��=FFM�5= (�      �'��P �     0&&�	�&L�&	���`LM&L�LM2100	F����L'���d� �h&�P�h��Y�IP����$�G�_`}߅���0�����D:	�0E��<�!�Y���\=4j\�����9�]x�-���W�
�
VbZ�������QC�AR�
 @ҡJ�-��qÄ��p�L�����b	�!�P�v�����r�����!-�痯���:`3����vӗ�5��ɧm�z�GG��	�(�&9lR�:�q���JS�����$QEN�Oi�(����	�:�F�����{���AeGC��Aq"X"�}BlC��!tQfL��"�c�RgLnU�2n�ش��J�1(Ջy"J�����CVT�Pxm#bX�1a�(HmQ1Y�s�]��4�gJ�I�*���:r���q�JU��N�D��a&�1
�V�l';��4U�-U�Y"��	3,)d�+W�#
�b�Q��0��`ȭ.7�i(å�M��l]SL���`ed[�����y�`��m���Am|�}D���|�W�g%����4�F2pcP:?�R5,����@�3�P]�*gu ��Y��a���Y��b�L������d�F=x���v���n����x@��'�Qw�	L�{���0�2�+����#���G��^�t���x�RR��?��뜭��*٪�&o�r����hlR7����|�k�Z(�=*W��'��G��&�NK��cd���A7r\X���V�ң+�$�'�{�y��b�v�3��h�(��w��K<q��{0]�9�P��_��{)��CT��t�Ri����fG�2�`D��Β��&kȿi�qzk���+��h-�%eE��E{ã���+n��L*��ީ�t�r��.@��d�� ��RN��G�
�y!�b��s�}K�6;$�o A]<Llc�/��>�~j�9z8WF;�ϥk����!�A��{ ��s6��-{=ȀDm ꋐ�x6�F3��M�Lhđ��w'CBj}��H� ʘR�=ЏR2�U^%A&�%�N��X@�B9��	�zj,E� ��� ��i�P��<����EA�����S�T�k��Zo�Z���c�'�Е�bytu!%��]A� !W��c���ߞ���E���f9*m�P#��2��7������\sᆞLf{h�=E���Z٫��s`,h,s��2` ���ݒ֍l�7 �:Z���A�vZ�1�B�@t�H���XR�䜴� a��|Y�/�)-je;��a������nU�1��9%��BG#M#=N�#�rE8P�2�0;