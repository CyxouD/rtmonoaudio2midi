BZh91AY&SY��,� �_�Px����߰����P�9�F⍵#Z�BI	���M�� �����i7������U? �J� &   LL 	L�D҆����44� 1 4�@sFLL LFi�#ɀF	I꞉�Ɇ)�� �4�4BJ�=�$��DBC�M g�;��|�����)2�\MC�n�1 ,0E�mCH���rfZ:����_{t�snL�ջmV�j<2�6oؖ���4����*[MڅUJ�P�c9���ꓚ�$e�a�x�V�ف��B�X�6 �.w9$$��r�.�{������&����xz�]A�G����c@�1����쇫I,ԴR��R�3����'-���WUKkLě$&�<1f[_� �H���Şl�F�e���Գ�ZikLa���hƢ�`R�
��А�0�D�_�j��Ј&���`��P�F
V8X
` ��R������Q�J�X�Wj�fU�pT ʨ�]�"HP�����"D��!UQU��Y��M��$͑��jTv�:�0���D��fGg�!��BL�҇K�(D��1���y9_��=&�T�7?G��$����$�@�"ɿ؟Y1ݾ;F*����(�nֺ:g"���2�,H@�)}�,�Fa8�	1t0�����baT�6Vw��g 0+�qV��ߌ��NT�vX��x��G���g�Yw�������yq��.�)�ι鶊`%����~e4i@����1,���xX<k..z��x�מ��8%�[�ä:j�a�!s�����	z@����MS���u�x"ĭ�'<~�.Ӳ(���ϝ}F9w =�� J_4���Q�^��FפY���.���e�k�S9�8	N	���O}���_�.���6P�W��|)��"TJ �@ٽ*��:_"ӂz �'dq��x�&���	�(O���A�a�����m%����X�ns�~$G�Dw��.�`�%)(d�}Bh�J9f���t��r\Lݎ��-CAc���1{rF���Yi�A� ��ja�a������{(D�uk�����K$#y���.�U�HF��c��B&�tEHh72�E�T%��1��#!4�%��j]��HD�e.w���n��.FQQ����c�d��c��.%
��T�ׁ��%�Y�
���@���������;�:>Ԟ��ع͞!�8�y��H�!�Y١*Ɍ�_.q�5�=�/v����������Of����l�b�CU�(Q��F��$�0o۾pOn�齆��8�J}
���j���t�%���H�`���v]4X#�1Ɓ�Ia�ghc�m1Ә��#Q��eU����W��9��F�%7#,�\H J�2?S%d���of:�	4��ϔ-�rE8P���,�