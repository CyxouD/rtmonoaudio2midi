BZh91AY&SY�X6 �߀Px����߰����P��7 �9*�E�(BI��$�E<�=OC('�2OQ����jO@
*  4     D!"�4�CC#��@I� 2=@s F	�0M`�L$E4�dL��������4 4��K?Ƕ��"��D! �}*�!.���Ꙇ�?bj~0T@�(����ki���L�GV�,%�U��K?0@S��Ӷ����ʕ��ydj�.	���MT����m���t�s�F�U2�1�{�u�Hǌ�o.�}u�ja[�(I*�@B�.�A��^�����$�0�����.g���*�7�l�c��v���9�v���:��!� hpD��'�z&x F	�f	Y:��@���W�b�B��G!�% �T���Xţ�Ү�6�+Í�#�cR�46Ȕ6G4�U�]�ؠR2�D�Y�9�2�������$�b�:���8k�D,���r���Q)�i��ƒZ���
��P�dc�XP��&�Fɪ��^	�ou�lj2��ma��)���?Z�v}������6�lBPA7����){}:l�U���#�x�L�nlk4� 7BP3���0� ���6�e�I��aE|]N�!ba`�֩�efL�&`,b�-k��{IF��xi�g�G��L%���?������~^�8��������,ڤ!/����̮z��PI���VSg�������r�b���ߕ��		n��8t�M��?�.qZ�t6n]~�5���j� ���/�NWq:d�تe�<����P���%g2\��p�:��R)�R��ӱA�g��K���wg`�������-��Q�b�UKP�%uٮ�iCD1 �`�H��N��L�w�;gG��}��+5"g�S����"kOb	�1?J�͠����*���!+�l9Ţz*#��[�HJe@q��P�3�N:�q���I��X�T�=K�Z��F&��t��h�7�3 BTKS�{�3���s���Er����7G�� �!.|�U����k�����*��DXCA��YJ��cE䍲��94�&�ߎ�"(Yd�8k��,��Y*OX�PEZ�f�t�	B�G=���]�Tf����u�A�=$��g���z��9�Ϲڕ�Ai{��_�h��#�r;OIպl)A��eg�~A�1p�;�H6�	9Q�K�;�H뺲�7QZ�,a�Յ7��JӚ�i�C�u�3՚�j-`�\�?X(�u��}J�:*����mW5"�J�-���V�D�r|G�9�*�7��V؎���RpfA"�F�����v��^���6��3RU9�l���A!+���b����s�gBFv�F��fPя�.�p�!԰l4