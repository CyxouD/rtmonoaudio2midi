BZh91AY&SY�� B߀Px���������P�q��uƙ�;��	$�&����<�C'��OHh�dd4�A����*�� `     $BOJ2Si!�<�L���A�6��hSU=�?T���������40M	$L��'��a ѓM��F��Ó\Q�,
�Q���)���S���{he� %�jU媇�Ȯ�	zE2@�fõ�W
���?���@S��+�w*�,�����JҜ�)��:�Su�F!��9p{ucsěj��6َ?�~�$f���W]Tio�A�a�ȁ'G3В*=�ܟ���$��:�)�y��¶7�ZM��0�u����,�s�-��p� �ĉ�`�{�2�j�����/��d��vj󅆌L%�姛%\۟i*3�a�.b�k!9�#��vs�w���@��dd@��%`�,�D�������Y�J�W$����LZn�,�t6�K�"ue;K��,�ֽ�M0JC��9, QD�J�Vc5TV'Ep����ԖV��3��$�^�A?�r��sZ��z��oq����{m���( �<�
{IK���º���2Y��cL���Ϻ&�E@(�� �<�j#�mKU�tA�t�-�-0�X�� Z�Y����O�Jzi�~{v˖s��6xK�ww�y�;^3������:1RI#��vz�ʳD1M#�(�7d�yv7DxѨ��ﯺ�Q�=��*.f5 -���ۃt���)�1�"��RS���h�ϡ�fN�Q�)���$��	��ӭy_��ۅ?4�(�Ks���s'N�^��mB��f���3�i�t��ݢY�[]��[g���g%ώ�B��Şd1X�;�#��O̚�� Н����"I!Ϡ��)�dT�R�s��a��a�������J*e��$����Ï�477���$�``��3��}ፕ6�a��!�@����.K��)�h,��N�|6c����tm4�$F�35�l�-�m��9��L���<3\�Z
�
��C�jO,�rl˩,���Z!���)��<F��rG���'s�	��_��0eJp��t�#p��[�+�)�2N�%�7k�4 +���@�Oe�ΒF��8=(��Ѡ�P�e�s�P{�k��
h ���9�{���hd����z�;K}Њ��a�&,.�8��T&���N��;{���������Uʖ�׹WleF[Ց�: �a����,��V�邞YDT��V�[!�A1I1�5�C$�5�������'�8�h+m�T��Ki)	�r6H������k� h�ˢ�p�l���:��~cJ [���-��r��g�&R9�i;Gg��.�p�!j"�Z