BZh91AY&SYEH� �߀Px����߰����P^8�DmΣ�M��	$�&��(f���=&F��  j����i2��� hh�  DI�M�A����F�=M M4��2b10d�2 h�00�M5 ��ڏHh4 h�MV
~�B�S������b��ߎ.�	:cH�0�� S11����L`d�w[��s6�]�޹XuAGN���Cƪ8-*�oȇ:f^�mm��u�i��P�����YA#b�s(W�x�P\*�r��� �f>`ݯ��uod`���o.m�<��}��2sV��f�x�^3zlo�L.&E���+�*hP��AQï)� �hhs��mL��w���J5��uʘ�[;�QFT�B���h@"2�jC�$�*�LB�$4:����p���!kJ)̍]�RiR�;H	�D�$a�PN%0�(��a�ZQ*^K��6�_Of����66�m���PA5�ҧR%.�
�*��E�,�3i������q(��R��ZS�Q$��@���/��� d��f�n�Y<3�h�d�7lAڔ�лo�q��s.��eA_����E���Ǉw��S��ۋ6U�HIwf������zIP�,��������QS�T�����"�c�$�Y�Y�7N� ����n�6$�P������}��]J]jg���Vs�G�tg�V9/�8���	)�E�m�}9ǁ��[ʘw�]"��ѱuF��1];n#ќK(཭3�_�?�SE)-Bx��m iC���`�M�iH4��5�7�bٓ�e9t"�5��c���VR���Ɔ��~+R���c�7l��
�-�vf�X�>9b�$����=gP�8��M�@m��zXTH6�)/!�q@ō���}k4�]LA%�a�a�{dxotDs���e�ǳ*�,��24	-�W8���5�s6L�"HڂY.R!����la�F/R�Lr�b�A�}��TL ���Y@�%m��9h��T@�j�Y���D���G�:��a��(�$�ZyI�yr�Z(e
��=>2�7H����pAYs��y����P��1���������h��+(=��k	�+F��k���/�]&m�1�fJ�Z��J�>pf�N�z�h|@2�1�,K����=�"TρEP+���j��\�$<��E�0��	(�\0�ZÓ�X4	���*�(��)	�pdA"j���ʰ�Q�\���i�o=�J�#�.'lJ�d{�Tgb_[�^�ks�8Y2F�ݶ��.�p� ��