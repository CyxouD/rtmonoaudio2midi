BZh91AY&SY,�}� B_�Px����߰����`_-����BI�dɡyMOxSj=CM�yF��i� �? R    h   ѓ �`A��2`�SĊ�i�A�� �� ѓ �`A��2`�DBjhd�S�2�Cj���!�@4��i����~Ԓ1"� J/H��(�?5�����Q�0lP5>2��<�$#�,��ń4�0���:�˛  _r��p��A3"��RH�ʲ��o�$@ �n`��P�8L�"d2�H����������J� ���^����z���%��^(4���� "�Ȑ�B�b�ۼ��$� f��*-��{=kN�x5�&uH8z+�v=�i鎣�U��[�w��*E/%FV�\�pК^A�Ͷ�H ���h�	Ӹ�h�׾�~��H�`�G�C�	;�2�%pj'I���V�$� �t�N@���Sd<�c��.�"����퐈QQ�q�{K�z��#���B�cz"^Z�ZB�a���E;:�U��"�t��X�T�	
Z*f���r�U�,
��a�Tl���SA�l0I��j�U��F��z�6�N7{����˖�[�2�l�;��<ηI���cx̘���TB��Ա����U���8|ÒI��km���Am���%/×���V{�,�g|Ej|�V`��,�S�w�4�8?xJX�i���b� b�¦�8�;��ɅɅ�W�S[ZM�d�L��~Q����Q����k�o["|��>6��S��������s���4`y�%���R֮�.\�+�B(�}W�O�rmY����5%/WQ��>�6T� �ggM[�t��pz\Q�u�6"7��OA���־dU,>���r�k�#�=z:3/��L�Ļ@A	rcn����Y�"�+Ӗ�PPd��{�G.BR�wU��Ｏ�V�#O��9��ɰ��1C@^4��1)�= H4�\$ʐS��(�0>�F�Ґ9ȷW2fxz��$F2��:�S|�%��YP^^  ���!�r#�H�u��L*�Cb���mj������)�xJ]9����05����*m���N��v�U�� A\��Ǫ_������eq����Y�`k�If�x�/X�:Y�q����P1X:��}E}UI���t��D�ND�wʯ�D����Jp��8U#!^��qU7M!�D�[�x� r��lA5�o�����լ��a+3B�����T��>.Ğ��k��FQ�4�L��B=�i��6+������L��v�k@@�>��9��Fڨ:�f��bT��*��1P �
T"��g�y����e������TX}��\��xXı�/e� ����f��ق�S�*�i,���V�1}D_y!�$O|l�诬�DP�v��A����֤�9,.���T3#��M5���sٍ.rF�G$xs�_���)�d�