BZh91AY&SY~�� �_�Px����߰����P\��{�;����7:�	$$�L&I?M�6��i�42dj22��   2@  %=D%<Ih �A�� F�E$G�#&���M ѐ  1 $P&����0�F�#   ,�Y�(N)5�I�,}����L�"&��*��1 �J)p�ch�a�Fk��m�޻���̤�I!f�im���:b�Y7��@���r�\�b�	�5���i%��v�/�
��"YJE	��6ӟ�}�U4�l<4w��y����i6��i�{������6��e=y�	,4W�6T��\ĳ*��|�6��:��r�����M);yZ��m�6�`�248��o|T��,Y�ÃR�z�гE���TUmg3�VBn{���  �D�"�
�kRȴi�qe�a;��vg:�j�3:9��N�����듛���(�ꪠ�IX��⸊���x/Z��3��ᙽ̘2W�3`8R��ߍ��ZgI��b0�$�L^&0��1�����Z�`h��2IPʆ)k:��(���<~˭�i�^���Ka,��(�������p��Vm��{B��I�)$�mXU���(�0 ˮ"cl�{hO�w�dG;��]�8��EL[8���)ǀp�`�	���wq�Rlhhز։��z������أ�tѫ^l�b���I)u%��֊Ƙ���F��M�O[��yBCܳI|�g;��JPN�Lb�Ω�b��$E�_	�98-������RSBA&�16���� P�G)i�d�")$�yL�L���r�s� �������X*خ�ir�U�T���H>�sճJ`��@9 ���i�SV�L|�%�P�Zo*�Oq�o�8�b��r#�޳=��Jw�1��D^���T�F޾I�^�m�e ��đ�$��W@A_%ǁ�q�$�h��A���+52:��dHdI:��D�}dDD�dʨ� g��4�HڋFL�2�,�TV"i7\��` &.�� �7-%��$�$���Pn�ұCQ�`������<濃������9��=���qorE����ygD�AZ��/�``�$;w��F����[���	_U~k��Z�!�:���1 ;W��7�����뺬/��AewLV���)��we��B��qyؒV���$�ǝ�$d�(�@�r(����3���B�" �H�f�5J��@�N6r*�b�EIȻ!�;�� #2:˔�b]���c��H��$i���?���)���0