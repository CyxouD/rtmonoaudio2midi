BZh91AY&SY��* �߀Px����߰����`�}�;� ��V�S��%BIh��L��i��i���OF����4  bh  sFLL LFi�#ɀF=BS�FM !� h  "�&I���@ �   $SI�����
i��i��   hF�^����H*�_�?�s��?������J�F��j�N����0E�80�H�
��η�4�$�6�Β�|gD%�SY��-M�0V]]p��@)"�I��%�yu)�*JC  �xfdD�@���ԙ��ad���0jd����/ے��@�dw�����'{�����HE�9$�����='Vꦁ	�4x�כ7��ڳU��LI�b�pr���lZy�sSR�e��Y�:�.A�k�<V�jWJ{)�kB�]��[ca%X��A �D�3�Ɔf��1G�fg�gj��o�\ꋀ�D��=jjm�B;�V���sx4����j4C�C��9�7��h=CV�*�麊2���`�p���$�S`.� MU��D�"T�p��n1#q�p<�}�\%V��*�"�����ޠ��,'^P�2.��4.��1g2X��td>k��C*V;��i���ZקgO1.U��MNa��0l���U|���z�ꥒ���g*Z�Nւ��B�"�&w�B�A2�ث�R�aI�<�k<�q�0�����x&b&t�è{���K$=��r�J�V͋2�Q��:�H 	0�'G��K��QT�/�s�a�ms���`�
�!��IHh4�ň�QI���yd�0���X�+q�ЕXD�G�kBC0�lM���vʞ�T�_�o�=뢓���%�ጳ����U�����I����u%�*Ĥ����?����������GƂ;��uDx�Fdޮ��ߐ�ȼ�<Bm�t�M,����H4�"G��"%��1|؏<-�	qq9Y�Ke��n��ѧ��W�c.tI.�T���b��z�4h��ᣵ�~��	�ۯF\L��-ڙ׿Z�Zkvo��kt�����,r�fd�I�I^4�jb�\�@4Zr'�"�����P�B!�"���L�b�&+ă@�(�o#���+(��B��� B����gtx��Y�BB�o 5��i�SV���s' ��L�.�9ʌ�����D�1y�^��`�%��e!Fx�fk^�O�0n1���c\���j��̤��G�m�R�ְ܍(��Ax{A܋�4HE�S#KlcE �DӡbBRp�w�$����i��9������q����hR�i�c�V��j��	�s�bF4Y�!i�R��V�����{?ҘuH��v$�-s�5�4�α2F1��Ύd��4O]���!� [�=����C�;<?��o��\f��`o��"�õc�B �5�᤺#-R`�Ұ���Z�*���lT[�^Z��6���X4T�"���;�e�U�8���Q*Ԁ�	�	X6[@�V-{H�j��E�R�ʕ'#&f��b�m�5u�ϓ\6o��5��9q�Я�.�p�!w�T