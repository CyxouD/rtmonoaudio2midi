BZh91AY&SYkcA %_�Px����߰����P���3x�Zd�E$����i�4ڦȞ�e<�F��F!��ѵ����'�  @  %4MAF�@2     UL� �  �   	�i�)�D�ؙ'���O(hhѨD=t!��	�$$�~e������U&X��EA!�a�/��S��U����4������=ف#t�+����@ze�#]F�p����(RH�J&)[8V++�T���G��>r�^"�j"�XCy�Y2A!��e5�ӽ�'��$�Y琄���pn�O���j`��0�||�ٳ���r�'���2�ٺ~:�v2*R�T�G�X��Q_�?[�rh����k�qM�p�B�q`l!�R2my��R�f�{;E��B�Q��K颻%.AFM�v@ �#c@�T:v�uzQ��)&�\#4�zj͹��f/L��W.%q1f�\��4����R�Ze�]�"b�0��*ԯK.�6S/wm|iU N� $��-~}_���r�BBK�$�@�fr*����C7.�j�$aw��N�P��p� �vtlBD8�w4����71��CF/����l"�I�}����h&��[����I(�V̸��:����0��2��w�+�_^����D�W����`�W�$v�����*�; Ne�*�G�����庒��2t-~�&So}��ː�±糤:b�yЉ��G��~u���>��
)J�Z� �����eLp�n�^c3I�%�	�Kk.�s35F�$SIs�}�$��j��8�+f���눵�Y|��v»���Ul�)t΁�!3��F "���:["��=�T'r87�)$	YJ��:f{�y���\��Q$ނ�dUS_?X$d)��vmD{�G���0hH��A�N�n�*��	���}���Ք��N�!�P��6���A��2S/Y��Ep5��Iccc�<�@{i!E��4�-��5d����	�Y˚��F/���r�L/h:"����ZH�����(ʢ-L�2h�������U��� ���T���5c�)Y)�"A��L��^¢!P#�`'��y��#�4j"�^lE���z|�����{�rn�5B	�l �[͜l9�6���7N}	F�0H{.���2n��4��T��U>�w�o^N��S*ҕ��h
1��ռ�&�?���o��+a�ؚ��4�6���4��s��H��"��8dc�`�
Vfʬ0�n@�C1w=d[i ��i�z��+�D�w�]U8 ς����	u���H�m�ULY.�Y�l�$fi�q�Ce�W�]��BA��8