BZh91AY&SY;�8� �߀px����߰����`}���JOt�W�5M�'��Bdba�C�=L�P�hѵ��) � 14  &��L� @     ��T�       EL�h h �   $�O&2�����I��z��F��*E3�=Tl�J�%En(,��c�?�յAd@'��0���)�	b0EX�70��Fk�ֹ�t�P
%P
�Ԣ]��D�i�͒MP�d
udń4��V�MB+	M���;N�&��I$n�.�v)n�[�rmq�߁�βR&3����Ӆ�0Hf;	���%ZZ��f���HB-]�f/nA�]�G˲逄��2o-7�d�u����nm#ZP����&R&��,M)9�N�6��Mc�|W���P���~�ڴʈ��u:`���N���`l���P�Hp�	�MQ��]t*M�B��pƯ3�",����%�h��9ݡU�32�$�m�	�{�)� $�Q��(�è��j��d�!�����jP�����H�D��'X����K�B�����B�]����F����|��I��U2$:����jc
��a�-��D�����Iz*J*l�9BY��Z������T�P���TgW$��S��V�U���\A*Ybī��HR-�b�D��[���9-^e�m�����h� ��HH[pL�x��ѓ�1�#w/)�-�T�`͠��(EIʑYr��jj(�U�MU=\ğ����H$�I$( �w������{��8�U�g�J�[U��З�IAU���F��%e�{�ET�@��H&��Y����T,�Xav��[#I$�2fO7��7��a{c��*��zV��b��\Wl��M����}�s�_5K�L�	�k�:�/=:����e�&a�$k�e|�Sïӂ����,׻���!;0�U��Ϙ6F�@�9v�@�hl/Hl�w}By����pkDҿ���C[���"<�E�_��1̀���(����"��3ZgQKY�F68����޶�eD��j;3��,w�5v�B���n����)�@�i�D���A@Hs�1�邡���'�QA�4��ev虦���#X�l��$��Į8*����,
n]���N.~��B��,���ک�:+ƫ��=�RK�������`!��b�%� ��4e��uLx���h2э�{$����,=������њe�T��$%�/V5�p�!�<�� r&�b.b�	p�1��#��Q;š	@����0C$��B:������i�h�5���Az,xJ�� v��l�&)E`!<+w��eE�C�uD||�8�[�uj�R�3�ۘfj�H�9��vt���	�z�#Rbp��<(Tx�۞''=1Z%�z62iA�6D�0o3��m���1vm�g�կ�A5���sV]*z�*sa��+�����<�kd)X�P�Ukו��xb��{�%�M"��c�.�e���i\�3�f����5#�����B�fG3�6$����.rC�2FY���g�]��B@�,��