BZh91AY&SYs�Ӡ B_�Px����߰����`_���	J^H&F�ML4�?L�T��O�H14��A�~�ID2	���44�20�jxJ���4�     9�&& &#4���d�#hɉ�	���0 �`�0�DГM��y����4�@��Q���ے���zWH)tJAb ����E���0���!E�@���B��a1	�E3��};�O���D��=n�C��\87�6jh�j����7�8���!6`_b8R�0�cj��BA$B�"� ��J�T�iUA;.��H���d�_�I;1�ۤ�U�\A�0ظ�lE(�t�� ��g�I���P](���>���		3ϧ��:s����~�?%��@�;�#���Ĺ��Ѯ!?�YUf`�tqŴ�r#�sA��X�"��D�%1Lq@�M()v�Q �n���&��8&�������)�t���(����p�Q�`s/%$_�ޗMmwՓ�K�\.���ͺnT��tyzm��jD2:��,�(�΅u�dO3h����£�ue� ���Cc��-kt�g`��A�!�kb�.9�<�W'N�LT�3��{����i/�&,�f�l�[	�f��g8h�����
b����R�73f2bT^��6I�0CjvL�c5D�+V'�h�R`�nT����lh�+!���X j�����%qz��t,�����j��bH�fA�e �����p�	}�T��A�x�UbjZmL�&��{��oXE����c�3:4�W�[V����/oW��NI$�TZ(�9���ŗ���d�|���-��1��D �_�V�B�B�ph�l�P7�E�تBU)��qE��#m��>v�́�r�p瀂fB(ʍk_��3��9Yg�~���t��7�O�R�/��������Y"�1��"���S�_���,��LY`�U��΢<v���<hУֻ<��û����iI����q�Cۤ��O�5�$^򐒗�A5�k|�w,����'<~g.G}H�
��z��a�П�HJ_�X�h�12uH���(.�qQ@`喵��S�v�e'���yL\%��K^Ѥ��2�C��@��-Ԁ�Q^`,��[��Z0-����m2#�[
,��~&�3���8Il��U�8��6j���(��q��W�+}��g��oG�e��T\apX<4(Qu`��H@n9�xL�zۛYY�A����5�bl��dڱ�=���20�0׽��|����]��|���L\���@���=�n�����t�R\6�$�*!��.�d�[�HB&v+qv`��@
���qa.24l�wR|�)��ݙ�d�;]��[Z�7�0*-9�-������^��!,���D�qѐ�P�
m�~?o���u�vEl���k����h���H�9��=��S� ���M�-(w���'@�ӗ^-���-�w��4�&�c
�b 8���ɜ� �5�i�#_\�-�<G�
S눫(>uT�T���h�Z��|�X(��/S�Wrn�6���*W]I��]��t�<$���EV���~U�v�H^��6�ݨ��j�#�Z�PJ/	�T��;�!��E�=5k)��Nһ8�~��H�
~zt 