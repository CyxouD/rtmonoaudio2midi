BZh91AY&SY0ay� O߀Px����߰����P�9n��("�P�$M����F�6��4������������	�* 4a  42� S%5��@=@�    ��b�LFCC �#	&"��SЦOS��hт�ɉ�Є�})!U�I$��	@��=�� _�����.`�"�	�aS���|Ē�`���ra"�.k��[��p�p�i<�Q��2T��L�U!�������q$M�n(���WZ�N+��!V# ��Ʒ.h1D>�$	V��$����Uyz��� LɁ�wzO�6Ӈ8tox�-qR�|���>�@M�-ׁ����U	�f�c0��J�
 Q��ٯ`�
Ʀ/6C�Έ C�C��|J�� �m0�H��"����+U�9��@�ґ,� �"��@�UR]VMJI�M⊇"�K`h��J�D ���
�ʆ[�,�u��"&��S#���ج�Ew�^0J����d�h��4҃AW7���K�EH���t����~�}�I�O���@�c&��<d�rن�n�N�"Q��P�Au\ ˩�CbFT��
b��f3� &.l*c�8�P��aR�
�:3$P�1KW�����Fi��q�^s�k���]�_��!O������<�/���	p��ϝD|j��x�'��a��s��7�uݿt����.I��gW�VN�P���� �|À�b&�`�tκv��56}KH�(��А��ZΙ��"u˯w��Ā�]� ��K�ΌG3&����r
	�n�:D�qEw�g}�D�"}4�4!}Sv�/%�6��Tj���S=����Xi#s���4�:R�N��"��-�;�2� D��Ez5&j��i�k��f1��ʑ$ޓ�^���� +�s;����֘4���A�L7*^��b����dO��$��.�k�)9�b�%2�`n �4�)Xf�Z����lc�'����Љ_��L.���r͍$��wyW 3�k}xW��0�|A�!��Q4]EBZ���i�4�J���	�~�̐���)' �L#}/�j�(�PD�	UD��v]�D�@��	���ԏ � �:	�j�P��%J���"r���(f�ݭ��8���H�:7M�%4`�ϡҘ�8���0�Z �^�4&7o&ɂrޮ;�P�%�y/S���Gx��D���>�l���05�;6��k~,l~�feq8�6�a���s 
� �����֔f�R�C�U�z.�,���xĀL��D�ԍ��8*W6�B�+^� �I\��Ѝ�N��T��zͪ�e��V���wH��$rR�U���w$S�	��