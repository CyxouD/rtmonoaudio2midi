BZh91AY&SY��� R_�Px����߰����P�ȧ7BX�H&@M
{I��G��ɑ�F�4�i�5O�I@44 4��@ !SMM46���F��h 4ѐsbh0�2d��`�i���!�H�4OT�'��L�2zOS 4z��>m䐮ĊI$�)	�J?gG� ��5&X��D�Pü�eQ��$�0D��:XCH�Z�ȹ:��I�`K9��!���:�iG~�Hl���9qS4�1zlM���:6�d����2���\,��Fg� �UB�V��A�.�� Js���(.�A����ΫS M�?�}4h�<1�`s�푋�kJ�F��m2��o�\V�8:�5H~[��Cj�y�L�K��i:���0X�l�)V��h�)�5!2�E����
F�iMo���v���t�,��#'bq��q-U*  �©�B"��G�(�a�	�(��[w���2�p�
#�p3��-!
<[e�r������-K6���[4:,8I�,�D�bv���HmEa̪���7+1界�e��'����������m��4�	��R�Y){ux찫OE�,㈵��t�AN%(��L$b����%�� &-��A����X�Z�}K�0B��bƿ�����NUUˣ-�j����d|��3��~o�8v�}3W2EZ�<�g;�`��~=��W^�LUP�i�Gewc���F���uX|���Z�`�YV]V��>��������������	�r���
ϑJ������n��Eޝ;����� 
]Iw1�`�-d���q4�T,���3�g�t��w��JpN�Y)=��[�#$�=�d�5���ڠ�4X4 �Х#H:�E*�� �:�56\L�H9pɚ���[�\�x2|̱$�2��MT��@"��C�ƈ�Ȏ�'�/3 UR��$X��y���Cqh!�0zZ+&�6���Ae�"k�����,��|n0 k��0�^�����ϧ�lj�+4�+�34�\`�κ@�����r�Pf=`�4��#+�4ƌ$�%'rrhI@��\4�"�e��T�9���qb�<",�	�HA7Q,�x.B�B���,�6l/FP��ܤ��Nb�CW�!���:Þf·fVIE�׹ͦ�v#0mT�Fr�6�%d���M`�i�p-z��|@	�;�}GW�=6�{4j�j���W�Xb 8s�9�# v15�N&�_vM��S�ꂔ�DT���:�%tu�$TPcM��@
� TZ>	�R�E�9>C�F�B���H_���Ә�K��E�Gi���zv�3�(t���ڊ-RSr0�թ���fGa����n]�\��,�#~�6�
�ܑN$k翀