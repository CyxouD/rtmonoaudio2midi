BZh91AY&SY��� �_�px���������Pm�n�Fh�և`I3I�~��CȆ�yC�b=	��h���`�PP      ��4�4��@ɧ� h� z�� �`�2��H���4ě�mQ�&�L5 h�	���:H'a"D��
��p���;W� �|*��`�#p �0��)/����ch�a&�V5��i�@\xؖ~~�!�u��u�YC�X�� �dٴ�x�5BFl�3c��y�#���MaN�?AGg	 �[�I��k��]�& 69?^t�n��ֱ�h���Jg����˜��d�ܦg�������'SX
IaM� �4�'�����mA`Ɩ�ds�[��*���AFLB����ʽ(HQں��_Ue�b�i:g2b�!��&��b�����d��U�4Ԫ�Pd�B��d*�Zl�Y3�� ���$f�/v��WJ���';��(����	30��6�W� �m���F�m�@A6۾��J^�N�U�Yሳ%�Q���5,"�Ia��T&���5Vj�\ imaU�:A}p�aq�,�������US���o�3�#=4�������i�w���1�xyp�tۻ��}Q0���d3��ѡD ��w���NR�8����b]W�锁��VW�u{I�ì]��"�үu��;n���S!� ���3:�kVio�,xQ*T}��7X9�k#�%Kg���|�lڀ�]� -����ܣ��R�6�E6
�,�Hp�]��K��t�j\����YtM|<�+쉫P�n:o3��4��EƐu(��4�t��a=d��o�����w�(4�� 1+١3E幙ױ#\>�r��s�^���^��9�E� ���R`�B�@.D��-�l�l���i�I��TD�Y�Σ\�W���3�8m�V{k�L�� �M,lc�q���(��ʘ]�f�y�/54�;@W5�4����9��$�����&�A����4Ɗ�,I�R.hH���+b@��ʙ)N����R3J��*��EHA5R�u;/YQ IP%�����YM� 5�=��=�1'$�](�6F�����TX����n���u�GC��ޕ�� }�qrL�!w]���� V�.:|�ĺ�t�Z�;�ɥ"[t�'@�����Q�y�v��6]��MZ��B6ָ�-��M��u .`-�x#%��d����}�x�e�w ��q"DՍm�pU��$��-�����17�Eї	�3��l��2�gb;�[c��"�L�������ܑN$!2�{�