BZh91AY&SY�vm �߀Px����߰����P�8� s�R"	J�	��FD�4ЙL)�5LM1�=G����55P @ d   ��D�=F�    �9�&& &#4���d�#I&�I����SS�=A���=G��WV~_*���QJQ��ak��>���hc@O5��0�Rc	�E1��|�g�����у��Kd��)�dSh�\Ŷ�tyd�dU$�J�ܶ :Re�h�9n?oJ�� ��oE(V�����ƥ
��j�K&bn�{�nK�J+l4���������̀,�����^x��VƆO7�h��4�pt�G|�'�HO"HL� ���c4L�fC�<��;��"��֋�AyD�"�A�x��X�YBuH��m��H�bJҶ�+z'Z�a�C���0�ظ�[�"�s3*�'�U��-"�Ș�)��N^qOy�4TU���ň	H��(�l�m�q;����0�';���rP�W)M3l�n*6͈,ȦG,8���X�N�PN�L͋�h@x���t����6`�}_�(�A � $BQ55�Ӊ�S��~��J�u�E����cqlDPHM[r
Z$�,"?ZB�2��\��u�F[��C�G�^�3�X�|���u�_�7޻d~�{_,<�
�_=__��7�&ZY���:�e�b�	y[����̥��$�(?6H}*#۾��7��?h-�|Oa�7�!k1�������M�Q��Ë!��
BJ|{�m=S���x�K��{V-Ɲ�Iْ=FV�׽{F5b��'�)y����+'Uޘ6�"�bz�+�$=�L�á��YD��6JV����������A&>�9!��D�Q��y`���h���K�Fj1	}S���6�/BX��c˽���&��Cqc�g�f����V�����J�7v-��nr�m遐$����	�uW����I駥���vg�d3��g�"l��C~0b�W�Ơ�M4!9-9���*�wu_\�!ͱ��T���=`o��:u=3�Z� Ԝ�.��Xrٞ.%��L�V�f[X�1��-��\ͳ(!���������4U��bա�=�"M¹�=��9z�O 	j,z� �ۜ�(m�7D?��t��9;Bz
9ͮ��0u-��9�'����]} �L-(zz�O����m����yv�q��Gz����"�$�Iñщ�� sf=�)c,I�ST�>0R�1B��Kt'��Cʌl�� ���6��T�][��Sl�7~����䭵�Ǆ�pn �U�j��/T���@����r�p*ʤ��_i��%c2>e�2bl���ps�5�d�l�pW���"�(H@;6��