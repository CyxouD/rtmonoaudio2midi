BZh91AY&SY�mr� �߀Px����߰����P��[p	�4�emeb	$!��h4�=F�&��i���22mA�x�z�    �   	�ɵ4��4=�=OP hQ�9�14L�2da0M4����$HL����F���4 2h  $��[���@$B@	?��]B����S0��G�HMC�
����1�s���s5ɩqyw��H[d���,�AN��ۅ͔eyU�M��cli��c�n�Ӟ7ڢFX���?N��!�bA�Ne����d;9 IM.ׂ@�����y�a!3�)�f�p�z�Zw>����`��֞��9iתf��7kþk����Ϋh�Ӎ�;̺��C<� f�3	Y'[2g�uO�;ә�kw��
��
Ť�Sq%��`]Ŵ0t�Y��QW���h��ETo�gZ,���_tRvn���&
tZ�e�X�`KL#VS�%�U8(USh�	:���TNea�r-�����bY2m�ȫ[��YRJm�O���{;X6AaL�v��;�?�W��ff�ߩ��`�B�	���N�J^�Y`���(�2Yɂgs���<��A���3�H���HmfR��	��(;�n����Fj�S8Z6,ř=]Q�j��Vy��a�qܶ�����;t��p���x��`6�������y'�DH[�����=�)!1<�ʯ@�|��x��rJ
����s��T�I�$,Kz���8]"�hhlH_�l�r�	�q�\\�Vگ4C�[qG��X��m��1�(X�
n��X�H�*d�Q��Z'�}uN��3�d����v��Q��<�YJ��݃>Z����F��i�gL�iC``i�`�H��N��&�AZ��;`�B��A�F�$',K�虥�y�[ȃA��=�&����\��!^S�6���".�vD��!=������>(�-�[-�!��󰬤���|E2X�Cذ8���e��HT���I�?�pz�D����s�n+H�FB8����˜
܋��cig�
G���E�TO�/$h);���j]̐���+)' �\%���ʓ�E�"JrL�u�'��.$�
��&�뤭D�`��l&A�N���q��>Ѡ:�i�;�)+s���n��E�1�Ga�shK�$'����L�אh�HP�_�1��Fڨ3Y�I�iP⡀� ��]����C��m6OU/�Y�[-��5[n��1%J[%U�/�xX�q����B�1�z�q�Dh�R�c�r�LmxWS5�� �P�id>
��Z51B�흜��ԦQr,�f���A$*Y��X����a��Ƨ9"�L��K����ܑN$;�\��