BZh91AY&SY+&� u_�Px����߰����`Ϟ&� wQEI�	��jzMS�L���	�M�5=4T��      �101��&4�H4� �    �101��&$D �h�SSd�h�z���<��#!���h����B�$@�8HJBH^���}�}�+*2��*�	�a��
G
 �`�1�oa"�/k�j��ՎI$��Ɲ�R/v�Z�hg��,�G��1M_�AC0&����XB�UE�L�;9�	��c`�� ��k��
rT�"���l��A#&�2d�l���4�^D�)߀ym��p�4�M����8��z�4p�4��@ݎL��t玎Ͱ{t�6:�>>)O��cHK���a�r@u
�P��"K?J�w�<c�ǌŅ�U��`!���@"��b�` 0 uV����n�}�#E����j�hײ�������3-;=��I`^�f�}��ME��[/!).N�p�[���Q���K:5��PK�'C�Y�,�*!�f�4�@�@d�m�׀��l;$�� �!��4�$��1���g���r�6�-���li3
�1��vʔ�n��Z��DFL"8kմ���:����_��\�.��ve�����z���p�|����N��#l�5�&�sJ��mm��;���4O��r�� 9� HJ������y�sqjZ.�glE�,눭D*2�� 0`�i1�lR�� f.[$	����H�"� ��0����ad��������f�hJ�*b�����a(�O9��w.;~�愱��+��z>X|���bZU�S��TJ�Qz�@/+v~��r�nB�4�����&ߖ�|��:j���S�o�r,f0
��ß?Hzo0��� ͡��\@�/�p�GKy��Z3"d��'<~�+x���T�v;W�1�$��r@(�%�cUc@���F��M����[�R��%�)A;����W.BΘ����r�v��3�H%��K%��`��#�	�+��):`�:⍦fEJ��H�Ao���.��F2��ybSz�Kc���� �p�#c�@v�G-)��{ӂ#�	#)������C���h��-��o?���3K9C�����j�f�fx��U����z��~@~��8v�7�ѡg���	x�v�|�p�ב���0�C�T\CA�J.��<CLh����v&� �	��]���W�N��K�T�z���T�4PD�e�Gr�,
�;���25�� ĀYo"���墆�U�0=��T�{zz
���廣�l:�H�!����͊�1�|�<����o��ϸ3�b�	�}�s��G)8�jU�TRVf	�b`;+��� f���c��R`�Vx�FYL*
��5ju�	] ��s*�m1HC$�ZiXdl�U��A�t,��E��ٱ�lJC� 89�$OX�\��m� _�u,�8ۨ��J�#�Z�P
�d|��b^w��c��Hœ$l�w���]��B@���L