BZh91AY&SYm�1 L_�Px����߰����P��.�H�Q*&�:��A��LMO�����i�A�L�M)=I���ژ�4 F %2(�I��@4 h&�s F	�0M`�L"I��eOiOOT���Ȧ�!?T�FA�Y��j���U
P�Z�r��~��v�E�$X4���B��H��*)�����r��H�g��bQ�c
U�m�L=��7Y�$$��Ȝ�4MU:r�-��9U�ۓ�T%=iE#n�lB|��0��56���ε�`6�5u1 �ᝅS�ysV޳�ד ����nߤ���K��R�3��`<�wL�lvd�S�-`�Y|�k���Z]c=0kĀJ$l���k-/$��Y�՜��D�C-Sj��rD!U�E�K�1!��1J�;�$�&��v8uJ\*�T�ppƔ,Y%-��{�JY%=Dcr�c-��<��=5�Kb)C��h6� �W��Afp�� 	��j�2R��"��FH{��^�p1,�`)���,��4^4�9}��n#y$$$�I$� C9��"|��z=[�E�)�o4J8�(�F"����B�E!#�F��0�.���(�]X��@Ł�o����FH��b����%Mu�d�>��u���	o��������Y���h&y���͗���Ф �O�~[�%�� �����@�uv���ꠀ�Z[��v�/t���Ì�����{,���Rb"H �E!%>~�5�Ɔ��zh�Q�T>19]�m�<GF��eԼ�2g@yN�.Զ1�cD���F��G|O[:�"�e��dg;��JPN㶚^���e.�I}/�_I���P�@�$@���6�`����s]F��X�&��fy4��o���J2ޘ�����/r	�1M��s�5�eԨP_���_���M�,|*a���Y�`�h\��EdTd�f2����@��Ŝ�~!���3�\��V��_NL�� Q�����������r�b�,�����$��.}k����p��M�ԗd�	zbTCQd���ڈ�&+Is0-�Ehco�%��^^&{���x�Vo(���� ����1}&M�[��k�ԝ ���R�^�$�0��!������#WS�+`���ٰti$�(�II�N[�B 3f}h�XZP����f N\t�$t���;�L���o%pl�C3@Ւ�j�9�=���a�\2`�D�f��K�P����&׷�� \Mj��@�0���.a�kQD�r}#���B��A�-Uͥe�`�
�a��5�t<;���A�g)�v�iqr���m�A�܀�<m��/F�Hv�)�1O.������H�
�#�