BZh91AY&SY��> �߀Px����߰����P8�t1֥�[4$�L�	���j��U2~��Cjd��z���T� $�       D"$������M�4h  4�ѓ �`A��2`�%bjOQ�S�=ODi��4���P�
l�@*���Qi����go���]@L@�i��,�u�!�-����K`_,ήl�p��>���.��{lxݸ݄�����fq���v-
nL��ͤ�-)l��s_ݗ9�i�P�ڢFX׭�:,��Fj� Ъ2���x��R�UU�J��πk���nὀ�``����۷�����?sI�h.L11�s���!��:I��*0�<��5�td�����S��7������+���hpjҊejc��;�K�K.J��Q��nfa�Yoޡ�b ɋ~�Fp4v�;�����J��s�И.��4�E�C�gሔ����9�1��C�8ҷm��R�$�uVՙ�m4ό4,�Pы��%3�[�bt��D�^p�m.�(��Sn!rcB�1Z�V�ah��J��BBl�P�.��[p�3y�s�:<�scllm�[m�	( ���S̉K��߲����#K7`L�u��㡕YJ� ��E8>P����#�A�Pa��0L1j�3����l͚6e9s'*S-y��x.���g�w��ϧ�������޴�yg�L�;$[�_B�$�o���ȥ�	$�(>��U��G��|G��i�q;��2�cjZ�7�So�6ySx�H
�(��{9�o�s�_�ϕ1*��s��r�N��:_�o�1�"~ ����ͳn��[Q~TÆ�/�)^5�`L-�W�K9�����)=��gӨ��<p��=���R�:�T-�	d���	�Ґiղ�:��p\�#���аҳR	'9���&oda�/\�\0�T��s�6b�V�E%��T#����*SM���"+Z���V��U��s���4��`���Ln}�f�Ag�D�1sj�j�-xF�`	(١�a����zi�#�_��4�Lj�c�3<Q ����%��sT�A����d� �ΥQL2&�אe�p�!A�~d*%�C{VP!�D�Y#!b�`��p�PD�u͏�.!%
 �nYLl�qg��It�	 �ݜ�P�o�}��y��9�Bz�s�n�#0~G��ES�m9�r��d +4o��²����h��{j}G�̖�he��4Y�ӹ��,��l1;~��"t́�Z[#-�`�l�>0R�1e��UV�.�aQB��mr�l	*���W���!��@�_}��0�]`��xHQ��h���$μ(�A�Y�	^��r6f4�|�Ex	�𸮅�}�5��J)�1Mv�� ��.�p�!�|