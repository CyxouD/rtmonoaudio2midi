BZh91AY&SY�S'6 l_�Px����߰����`n��v�;�b���J@�AO$�S�'�l��i��0��A��JH���hd���`hEC���������F10� �������# ��M�	���dɓ#	�i�F& �"�����6������ ���
vh D�H��$�I��)��~��@����S0��F j0��]�$�Z0D��7��H�
��ػ�p�4��)��@�v͗��ˉ��t�8�,L�6��:����e�R���SSG*�u���cu�*�X���S�qi�(e���Ʈ�S0ރM��	I�����@�?���M2��w���N��v��S��Ě7V�����l�鍕iF�3��E���I��{bvS�fp�W!�`:w*fR���r�1�GNdJ��p�cF�L�ja(�w�1�dY��u���&.�8�v(a �HR�9)��fd�0�.\�j�J@�-(*�JY�ކKf1f������s�;���	��8j�e��E+�V`�m�'G't&$�+["�8B�0�=Λke������d�7���S
�*�'�y0kYOS3����PD�^��H[	}�V��M�t3"yL`���e���&�*%W"YG��"m�0͍��C���D7������llm�m��1!
�k�����>^��-zߓ&S8$�ņ���h�(4ZEDdPa�Q��5�J4���@����e�7:�1A\�mKz��16��s/w�X���Lm�_��CY�F�󐃋� �E_�UzO�������<�"��ߥT�f+���8�B)A����ۀ�5���<hУ֬=i��2�c@���Y�Ro��.�5�6��໼�w��ӵr`�%g�B$y ����Gq	S�5/������Y�@��r^VsbF6�4i�D�
+��V�P�0\�_6s��ħ��O}J��y�b��gœ������Z;,�M HM�(v��t-�p&V�����HiI��@�q<�&c�����N�_,"�����)��o,%�pkҋ������˕00�zpl�&��fX3h�)����B`�Y5�&�&���/��X��x����367�����ϫ�d���6�,����(qڷ����m:ާ"��{� �e"�]%"���H�l�x+F$"	��cQB,.f�8�ݺF��Ya˪�YBPB�R��x^c B)5p�'���"2�A�}�u��q
�����:�_�u��(cs�>=���Z���tyҤX� z-��L���k�@�
[g��������+V	\U�Le@8u�.!t����Q��`�y�v�JwDU#)^��U_���f��<�@�Ɓ��U$��ܦ���QE��`e�e�A
�"y���!F�r���l1�nrvi0X���e�i���#�ʣ&'���f6��2E���bЮK�.�p�!\�Nl