BZh91AY&SY�<� 
N߀Px����߰����`	�{Á �u{�A
��	��6�eOS)�~T���BQ�hh0B*~EU!��00L��#�lI�M �      Jz�&J�       �=F41bd�##F�L�@D�MLT�ꞣ�OhLЌ�F�}�Q���AQ���	@"� ������������$�DF5ׂ�C���8H�|
�gH���_U�B�Q�C���8 �ۓG�	�$���A�bEQUQXEUDU!�AU�UUAXFNig��d�kkV�"�¨��+(�#��P�n�N)<6*PK
3�f3�(&��"�31���ۀ�.Ѡ��[�����>}���ш��;�}m� �M��8�Ȕ���_Xʋ�A
�����!a^���ji�k�ʣ�Q���2jl^Tۺȶ�aܜwJV�Pt����q�D���|G��y�M��.Fݛ�۵��r���"�c���\cSw��w�/$�ƀ�)K���nVo�	-��f6��l�1�.�;Ы���1�o�5�4��SI��i��nف�j�-��-��.��ն��֘�R���a+,�e*�l�Q��u2ٺY��[o�N2�7s\�L�JܘX���;8ڷK���5�����1K��i��5;�PpC���kJ��u-{\��\��A��%t�1��:"c'�N�AE�ky�O���'�ox��Σ8޴�غ4��/aZ�����ȸ]28$�%'W���'#h�ƌ=��"��W��>35ԆQ:�Ίjb�L��z 9�V��k��8r��i�ri�d
��n&Z+��'-���1N��z5m��3љ�-�`����c�p��L\�z���8$q��7t fd�ơ��e�i�tp{oj	�����1Sw��:�6��+q�=�.k8)��������"��+��˒z�u�8pĕG4�N����q�`(g)�{�{�Po�L�\6UZ���h��לuD��X[m��dB����!,R �2j
�/.�7]�����+���ACI�KR�܋c�rq�^��5�u*S"rU�����ix]�#�4%��U�N��%<	��_V�~=?�'��*(�UPH��J_���Ė_��'����b�ۂ��h�tP�4�QBY�b	�1�
	bOt�h! ;j���_�n�?э���G����B�%[�ca���r�'*��QЮ�����D������I:&�L@p\__%dn<d�F!B���Ȫ�D�*\T�������������Y[֕yq��	���,V����|��>×h���"#� ����fӲr�?.����9�1r���4|�FWp�E�׹�B���f>;�%̝.���(�'�>�'�e5��g;�h����d���OYo\�%a�r�P��Q@䖍�� *��E�F_-,kz/�Fa2�;��i�(�n#>�o�K�r�ނ�%_8���+�IEx�B�#�3�-���wT��$��Bޜ#֥	��FJ���㬇9����`�k�yQ�-]�M��@p��W�^��B�^,36m���G>�_Tj�c,L�`����-�Bw��GD:�>��-Ipԝ!2L�,8�NE�B0����0[d�6����\dhٔ��sd��ѻ1U���E\(�mZ��3� �}��3�^�$�"#�}d�}�j.4�~������a�3��ث ��9�q�9���)��#������](�)�����lB���C�<>D�YQFq�^�95��R�Z��b)8v�E�"�����il5FY�`�d�?H)O8�����RWF�)	�(7�kf�����߁R�j��M�Q��3w�\�5�Sd:sI���,,�+Na�{jg ύۉ\��r2�ݹ��!
�dy(ɉ�8�{1��$md���8_���)�Q�H(