BZh91AY&SY�@` C߀px����߰����`?v���UT�	IBI&��2A�Ѣbm&��&��L�����De�   �  0&&�	�&L�&	������� �F��m@��  ���&L�20�&�db``(M54F&&����<�&�F�4���Ca��
�0R���E3J>G�������m`H	ި��%�A�Y4 %�"v��R�2�������ܨ�w�G��`m�`��"�J��c�H���,��(5D�m�DA�B�����b	~H{8A��� ��.�8"w�ƺ�n���܆༴���UD]���8���=5�2H``�_�F|��=�{x4[I�� .�����n�MZ�N��
�'o�"΋a�_�^"D���$m�@�a�@����H`Ϻ�a���Bل�Jݰ�6̱�w��������B-WB�����aq�)�(�Z9[kM�����D��	�1�D[N��+�ΖEJe�r��j�n�C��5.r�,6n������%���]�L�l�\�@���F��S �M5�EN��l S>f�����)�UJK,U�`��Z1<�V6E3�v;����f����Ӫ������cYy�A��M�����a�$�A'$�@ \a�#���t��*�dZ�Ȭ��8Ј2� ����Zb(A=��
c@�Jb�{�b��jc��ve.�kg`@3%KR�Mo��Q��0����pk:�D7xم���yO�τ�������?i�簫�~mNj�������gC=!S\�_�s�����T�ƒ����+>��1p0���pvA��r�� �đP;� Q�z�m<����j�\�m�����͐G�s每5��1�B�;�@C䗓TK�K���k�����6)Z>�f��������uBI:�8��aaRI+'!���X�{��*°�
҇X�a�M-B�:/�8��	�U��_���f=���CR�=ҺD�aA5����������	��\���b� B�mP�y�3N������[�ɪ䤈/fLz
cް�%4V��K�*VC-��3	@�g$$!7�u�'n+����L���6:�3<0Q:������8hvN�Z%�Bu��1i��Xr����0��JjY�+�Jk��R�X`dՔ~4N��rl�)��*Х��nҰ䘾��QŸW�� [7%E�2H;s]��'�}7��}cHm����Jd��Z�5��^3*���#i�{�N5�T	ϧN+(>NxN�@�62Lv�!ut2薅jT�ȧ��IÜ�b����5F�%ϲX�"�MѨ�z�uJ)�I#4�(.+x��:��.�E@�o-�%9suMaF��7��uٖa��='1L�*�����Nm�pU+��1>պ�p-U�&�AE��a�;��� �H����2����C�*�Nx�:v�ϼ4��ܑN$%�