BZh91AY&SYϹF (߀Px����߰����`\��# �ƪƌ�$��h'�OD�=G�6����L��Pj���� �  4  0&&�	�&L�&	������=!F��h�C@ i���	���dɓ#	�i�F& �"��ғ�a5Oԟ�?J0� ��hX���&$X��`IM	Ns޿� tt�rVfl] ��?�2@"�Q���4�0���ˇ�M�H�U8�"ϗ������t��<��frs�HM���*�,��R(!�2]՝��ǔ�v3?{,n���V(f�u6��Ŧ����32'�Zx �(��$	�V���Oq��ri 68|�n��>��m�*�A�a;/s��&��V�'ry�=��:Ʃ���LX��5zZ͢4��X��2b�P\��a�v������d�3--ylf����*��a�t��h�,�uB�R�ͬ��&�bK���il4r)�$�idw��+T��HJ�v\���(�TNQŴJ{� Y}�M���P�ivV�0��p�-�04�-�X�|0�U�M�R�8��ZZ�I�t��Ļ���-anLj�U98���:m���K�\����r�M���b�4�]-ͣ���9D�:�z�^O0�D@����`�V^�^������׮�2��%�l"1Qt;S A�ƛl�D�ֳ���ɨ�6���� ���#^�N�AY�S��e��Ēmb��C�u}da<�ra���[ o��"�/�'�/����*'����z�@���y���h i�T�8`%ף��Q�KAC�nz;O_�����+��7�r�Q��hm �7��'�q��o�����Zܪ<~'*���#�:XY��ҿ�s�8��o�@��ٛ�������}�R|��4J�
�o�i�˼J2'j�{�T�V�B�VNC`�%�l�� �遁�		���k�-pC �
`�e���� G�t�i��SJ� �c)op�oIb��QIx�H�y�do��D!Zp֘0@F*̈mR�i�Sf����$�=,t�bc%�H��%3T��NyҬ����$<<�lc�/y�|��&B7�|�k�3���%�j�bnbpH��vT�����q�$0sEH4B(����4ƊD�D��X`�j���(E�e�*N=�H��n]Vue	A
�JgY��@ "�C��POg�4jHb@z�A���)r���c@n����'����nku��R��1F�ׂU�@u�9�E�]��H=� AO�H��Ev�cѯ�촥�t�i	��7��Ja	y��t����0�u؟	*ݾb���犢�+��H�7��T�/i S�2,����HE�]xg��=�.��TI�l���R��Ij읜�EW�*PQr2X_{�������E,�����js�/d�*�k0_�w$S�	��a 