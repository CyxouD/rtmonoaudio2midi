BZh91AY&SY�� �߀Px����߰����P�9��8�*�a5��HC@����z����z��4�6��Sh&%4�=       "���F&O)�@� 40&&�	�&L�&	���J @�&�=OSOD�	�2 L�A\�"��R�E("�g���=�ޛ�!|	;U���)C��@�@K�"s@�R�G�����ˡQ��yg��}���>B���QƳC=	g�z��,��Az�E�*�f���5����+T��C9���ތ�E0܆+��vG�"V��+}�*�:�0k���u�`�FBH����]Yv��d�ߓE�������ٱ��7>xʥl�Z <�@u����L����My	 � �d!sB� ��{�&�G{	�yL\j���V"��iKa2��p$9l���)1���d�L���aW.)D�e�R^�*�k7 YsJ�*jņu-r��QE��HI��.�j,[�a�4Л�i3vI�ZZ�J��@�E�[�9ժ���z�{l�iG̨F; �����/�A�i��X�l�Yic���u�t������m��0�+M�^������׭`�g�����P8�A�)����bV��F$�y�ޝ�)#d\�<��~�9 ^@�6��o]��5�xFn�3QGV���u�����o�vx�������|~^~2���'��ҭ�d����}|�/)�P��s���RN[~��JJ^����S5��@K~U�=�?���x�H��� Q���⚸�"	G�|`�̬�q�������}�5ր��֨߱~��x4����U-�5x�8�2������w��%'p�i��¨�+�i����Ni}���iF�A���Ъ��
��l�f��*q�奴���b��Xc������!�_�e��&є�.F�ǳb����3�,���k�R``{Ӄx���Q�]j]{r�C�)�aj���V����IL�,npݜ֮����$�%6��0�=�>���r|��$�=Lg�I�^�m��Y���ڒn+�����q9f�Z%���!-K�D7J��6ݒ�uJbXˊ�����TK ��S��tF��2��x�u��	`�`�3Y�� -B�k��|�ʹ�Tw�|��{���
�S�@��}�Hv����PAQs����1�<nM҉�8NM�`�d"�;���p����n��I	�N2�S�Л�-��J�R"���f�'���H�@sXxdc�2,cό��A2��t�F�2�u+]8Dy)����!E�F[��(x^z��#`�#��h?
��dxL��B	�6���U-70���C9|��&�EN�k���px��fG��I3��cٍ�rF�L��N����.�p� $���