BZh91AY&SY���b $_�Px����߰����P�8�i���m�f	$�S�h�OQ���C�Hz�I���4 B�P=OP  i� S$iM�=@d�M?T   �101��&$H �j����4S�SAOj��ړC@4f����
}פ
F � rI)�B��'x�ϋ��#��UI�0lPHjz�󘄯"�mXCH�Z�ܸy}W�	�[���0�� �e9XU��1�^�F2���9���H[/_��?\�%:ت��v�>d�<�lC7Ŵ�:���r�oZԪHU�R���^u��{mL�����w�\;���;\iA�(ͬ�m�n�,�Ju&V����<�ؖ�ً&X�;��֬6yP	T��� ���"�J�����j�&$a,ɮ�`P�3�T�R���8����Gu4�i�
-����gv
�R\$���b7U2���.�&ir�ht�iB�0�gHm��k{:b%:0��%�U��cR�Y�o�j֩��e�0��tHTV�a�U0�����z�����6�l �U��KȒ^�g}���Dh��b�T�H\�֊ �1U���E66P�_!aH�$1qaS8��4¹����S�2��4=���6�ȶY��d���j�)����v"�ׇ'͗��w��w�cΩJ}X9������y��QdP���	;�#�G�؏4=f��Oq�)�r�b�$cX�ٴ6��p�9u�`���	C�39y�	�:��tjX�D�G������G��e������ 6����D��x1w=cD���Fg�F�=k��$�,�-�����	Sv�2�e�����9^���!��t{��p(���*�+_T6Y�� ��ˌ�(RH�يf7w�$F2����k	�'��P^[#=+=�p���$sbL	���A�J�tיW��&>�d�-	%�A0-V�`1�n�%�1�4s�|
U���%fP)n�61�'�>z��P�]㺗��Ν�f��`���o�_hB6>ϭ�0�{���k�M�P���4Y"2&�I\�%j^�1$"`2��$��B]TH�V��^�R�P�1N#���	������r���RaE���4j%A��J�0��!���5�����ho(�ї���4�d#����J�1�C�����7߸2�D.��Y;_�5��l��թP�VXb 8v�m$"�3T=}���=qс����b��pV2�4R[�m�]�^�"�	�L�{.X�B��G2�t[pY�6;�9�H,q4��>|���O���+�vr�^IR�L�d���t�H̍�EX���=��s�.d���O�rE8P����b