BZh91AY&SY* �  �߀Px����߰����P��n�#VZ��EBI�z&�I�S(��&�m h�ɐjziT�(��1ꌘ�#j 0������F� �hh   ��A�ɓ&F�L�LE&��i�i0��P<Sj � A�"}�"� I�B��$����~Jٛ���j0�>̹Š�M��{4���[�.瓚ے�*{3�ϼ [�����-]vt��Q}��/44�cm����އ')�W4����s2��c��ݰ"1���>�U�u�A�|�9�*	��wud� ��M㛾y2o==�W+����l�V���͎����A�������Uy�i`6�����*��!{Ge�,�2���-*����3��,�&���4<-�oR��U����!���`�T0k��ˣb�B�򖹃i&��.�C��2(`�*
� @�H����P�%�(d��'wT����@��`��
ʛM����}�x�	��m���B���*򔗟�����]�2e3�Lb�����5J0d6�l�T>F*�-ja ]�ZÍ��r-Xf0ѬxKX���2
�T�moc���Q���oٰ�^���o_��q�Ww��.c�wq���W��!aW��U$��ˏ蝖��&���'Aؔ����x�VV��a���u��f\�n��߼?�P/hm ?Plg-{�՚�.��b ���/�G-����v%DlяZ���y�=;�3�UÑ{P�b�-z��eI���9�8	J	ګ�^���a.�J7�WM@o.+�g�����Y�%��*��O�Fۅ��<mGd�}�0b��g�S��ŗ�,W� �a���C���)��J���H	q}"��$7O>�����@6�X*����T�˓[*Fۈ��i�b�H�X30��p(5���mu�ƹ��$�4	*eccH��n`|dB6r�+iŚ�+�@��-�{¸��gkS��΢,5<#24�ŋL,�4ƌ蛥��[�j�Y��`3EI�g�%��F�h�f�r�%�+%)�+yH�h�Dd�Yj/�$���E�w��M��U	:]Ȟ��k\��n��0ܲ�����w�^�J����ԄmL����B�li �F�_I��Gs/`�D��RWh���P!��T�w�&d�5a�
c;*U�T�a��'<j����	��5Ys�@Q���<�+�{ �Y��M_~*X�fwk��(<"��9�k�z*�}$HZ�f�A�m�Hب��0�i� �T.G��J�S痦-�a���#5n�hO�.�p� TL 