BZh91AY&SY�� �_�Px����߰����`�� �b�XH��I
i�BM���24�!O(�)�F��2���%@ 2h � �M  9�&& &#4���d�#jD�� ���4    9�&& &#4���d�#RѦ�T�F���hi�2z���4�&����"�`R�A��ŗ����OOά�@%�@yN?�<�8�	X"�P�`/��>��<rj�</�(Kd��ԫ@�����n.���F[��b���ܒS�L���q��h�G*��^0��ΩG b��|�(����!�V/ABլ� �?^!ν��ϲ�
�~��ѣ����h�k�A���si����k�OQn�w�^C�㰷xN	B�D̈�&��(�����b{��OA�%d�H�C� ��I�+ps>f�����U��{RF"w� �!7F�;c���Xsә7;OeqS/�Y8�I=�Uɰ���i�鹷�yS=u9�lz�Wq@���+\�(#�f�0�ח�uv��6�0v�	C��P��C]f�@i� �}�W�3�sI�Z����ZC0fL�t%j��Ι5q��[FMA&� ��vX]�\�3X�����{	�V�I�Rc��z�E��ԕbM۩lmɊc�����Y/A��v�8�J��*[9b�����Y� @t� ���^�;�Kǻ�JuJ7;��1��)	V7�*9	R%(�BhBHC�6�yD&� �)XQ {�.j��I�N�0�c������湋�/���?�ҝ�X��{�\�o8����.���b�?��ˊ�24��l���E`��,4�zzɕ$!�P�-��ʲ[�}�ȁ�qt)�S�3�݇T�J�mz-��<-�z{R�� Q<� ���x����Y�$��Ofu�n���^My�?h��D���Aը�C*����B�u�Q"f�{�Y�~�+*O���"�}��6���f��pѹ^��8Cm@���j�۔ᒀdҕ�]S�s9X4��rӢ�C�
$����5�-�5��2 ����JlFf%q�գ��(�6w.)/)��m^[�TI͐z���Nu��HP�^��	��%��z8��H���08�e��]	�s���k8����DFXmG���CŻ�J�v�������@��oܻ �����:[SC������D�d�*E�թM�0B^d��b����?}�&% ��ؐA�$��Mv��X3��Ȕ�D��pm�>Ң�I�%��X���6'@�t�Ӵ��12
�U]� �~�~����5�?
��b�����`ڳ2G�tx�T�0��,��ؘ����s�PmBW�\Vx��υ���غC��a�P	巑LT��~�3�������6�,A���]M��q�Tĩ�FQ���N��[����&�$k"���/��ǎ�6q찀�ʒ+�l��0�)ֽ�����Đ��6o$ߙǌ��j"�8��Şx�c��#;&H�x�yB����)��l��