BZh91AY&SY�=� _�Px����߰����`�&� N*��ٕT$�S�F�jOhd��L���2F�i��S�4
J�0�2b44�h1 sFLL LFi�#ɀF1!�I���6� OSѓL�ѓ �`A��2`�%�!(�a=OSԞ��~���i�@�F� ��Bh)p �GA�TZx����~�k H	��F�=��P|.A�	hH��R)hǳ���n�b���_�dx ��3��i�o��8Hdn���\��s&h�R�6� %�pL�6��]���()�[._�6<��/L-�v۶�G<�T����i]ƺ����оc**���P@�}y��ܽ��X���>T���rˉ_���hcA�`߿[_����3%��������6���,��c�2�p��+���� ����t�<5�X�a�:^���C����i�,M':O#�����ѝ�u��D��Q�p0WLK,ݴ���Asw�Z��]^P#*9u-s��ؗ""���L,}E�8m�6�X"�"(@3��V=-n5�nb.��pl��c�Νp/��js��$�^N��h� m6-�fe	�6en^�5H8�=1̛�L�0}�$�j�Hs2�u�H��4��Fr��Jb�I4�B�"���z�2��:b�gCR���U��s�s��X؈�����hr�0�rI��m�x����?����bHHI>�$�J+m�m}eW���{�׼�T�Fd�A&�$���� �AF�  z ����� ���
)�hr�L6Q�c�9�tDI�J�ou=��A9SO�>j�ͫ�Y����Ϗ��ww^�dVU�NW�$c�R�BGexyxx�`$�)�~J b��G�_�tG�������;����c@$�U�״6ɻCԣ�&!�$�)�Q	(�;�jvO���y�%�GBs��9W�{�����/��1u��>���u��	ש.6F�O%T�n����eMT�|�nr�ϜD]0�`���0]�a��X�C
߶�1�����+ 2"R�8�P����iu�P�K�O9�٩y��)J�[�s�v�^�6����Y7��&�χ%ȿ��<�i����X�����:�KY�v����[t��万4��]Q0\��
��q���n�Ʋ�=���HH�V��0�=��=�nh�}�F�}0�4a����#֢�����'<��7��.��%�R!��a���ۈ�&)���� �5���TK���-Y@��@ؤ@�E�1b��a�A�#�g $�)b�`�?2�fHH�!"���<-+0�Z���'Ps���u�TX�6�6��b�)�Q;�9��\+���> �XVPx��pN���j��|:5���u_��t�]�|!p�3`F �6C�y�c<&�V��:��<",�
�~��c׈`T��]�ǂ�eR����������!�A�bU�T�3�K\:s���KjN�cH?&�%��w3��PM�:�lp:����Z�p�����2b}��{1��#�1M������w$S�	
�3ؐ