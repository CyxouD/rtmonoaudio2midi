BZh91AY&SY�o	 ߀Px���������`	�/ݼ    \�6dūZBI	��mM2OD�22m b ѐj��*�   �   sbh0�2d��`�i���!�i�T�2d�z�h�@� 0��"Rɪ~��OBa=!������m$OҍM��4 1 4 � �f� �R�@���PY�{_�*���ָ]@O�*����t��֢�-���"���-�N�uZ��[^��!�~\8 �٤����VMo8�5�wf�ˉ��aA�:�0Qr�6*dNأ�vL'�āƁ��	�Q�"*D�A$���,�Z�lŤ��l�!e��2�����U(��G��+��k�� �
YV�����Ӌ<�C49�hk֫L���]�� ]�Ԣ!��p��n��EV@����ώ����[�9�5ӭIp�y���I�O^�1.�j-%�dL�T���>��7��o$�sn$5��֚f�E��{0&��Y�� ����6ijhX��,�����%�-J���T6e�0�=�0���/b�r5�ja�۪��`����*Lɨ�� |����Eps;Z YiSh,��G>�ZΖ�R l"|�0���>��B8�8��䰅r����&��LE)	�� �F�!��-�+�<���4>j��L π���>^�DC�H��d<aI[~Mj�lC���8�A󒺧�� �m�j��#�a{ŤY1z�
hҭ6�����%���B65�"�ͺW���i_p�7v�T*��w���\������g�-<c��pTP�S��	��":�c���!j����k�9�gC4p- �=f�H0�Jc��Z�-'G�7s6Wh����#D�u]��z�����9i�K��F��Ѭ��|�ᩥ�v;�.+�_a�:�sXt�x�F��w��I���uS�#�Ţ��r�	���������W9W�*��'�]lSR��@^A@��Td��Յ���92"7���n�I�����P"�LAA����s��MDVV�����U�=!B� �yv�_;U8:f��F%�F�sA�XfN��rޢ���b�����jå13����y�xVd86���1.!����
�B�7ohux6�^`��]��q��d�j���,��V\�w:��.�MĞ.y؂UKa#���X��:#3C7p����Q�|�~�;�Oa���v�L]���4�~�m�W���;8�������~a�I(  $*�����z�T�R����b�׉�S)�R^� ��a��l (4��E�"�gA��i�aƪ\��^�8��˻�o�q4l��p��<1�;)Ӛ�5�a�N�\��.��y!<;`W�����;�ݞ2.,�S���6өM	$��k���U��$�b�-�{�Q����@񨬭����S���嬹��$�Y�n+���7�y�]"�qđ_�$J<�c19e||��Ib��m��\���G��Fݹ�����P\���J}�ocF�����/H���i@`{�jWƦs��	N	ދ%'��d��K'�(d�4wB�; �#GQ�M$'`
��7-p�PK0NB�f%�[#R*���ra����N�:���l�L���/mk�U���8wƟ��u�x6�R� �I%�����>�k�u���C�i�_Y0[�����B'������P*��ݧE��*�gۄ�&����	�aJ������eP^w�(}]���2�nMX��E�X�A�"4������cFTM'��؄�z�С�0�8�Dp]#1aYd��R�:*��Jf���Z
�F�B�����LM	����*���]LB��W�@ytyN�陯{���l�9ͣG���<.�Sp�u�W�T"*�{H������I9m�,�#��OE��o�EJ���c,�$۽�^�,V�/��W�v)OU��|���a0�QU6�P�Nh����if�ܓ(Q��p���e�5�M�6qӘ�NF�	�l�%�\\d��u����ڤ��_���I%`̎��D��~M��J�Sz1Ni͠0���"�(H~��� 