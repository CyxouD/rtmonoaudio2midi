BZh91AY&SY{ӈC �_�Px����߰����`��q
 �u�!$B����4��I�=52  S �{#AJ��#F1 4a��"%�     ��'�􌁣�ɡ�    �2b`b0#L1&L0H�M!)�z������4���j���z�$/P��H� B�	�>R%g����$��,��0ld�P�����f6���*��}<�ӂ�I `���A�ێZ=#�Ƣ��eC��UK,F"cb�e�?#;��T�ptޭ@)�	e5Q�� �EMU�%m+7b��EDD��G?���x�	�Sq�Pf�׭�=,��FjdC�Vza^�����Z�eH�/� �n��Ϧ餀;{Rא\�H�o����H���R"�H�@��4�@hMI�q��C!<1�Y�����ijG��'V�ev�P�m�-K{���yLks4�Y1HT#Ma2j'��cq��,ݾꄖȀ+�iF������0����98ڮ��������;�%�,���!/2����5d�r/
�4[]��Vh��N��T����vunW:p霮JD��c�pn]�Ed�ĵUCk�6��c1S3��WRb�ekH��-A�	�CfUg�ckR�-��Xj�����Θ�MeD.0D ��M�>+��O3ȧ��E�(���$��{��V���8�3]\�''��������nԍ�̣�\T�TU�N�nw^����mAgDK$/D��uS�TE��Ͱai�<�X�4K�%�f~W�?+Ca��f\ٸ��\����5��+��NC٨B���Զ\�J� جM����b5lj��[t�7�		KJ�>�ߓ̹� @z@�n�e=���{j��g�"̖u�VŒЗ����c]m�� ���N`�2�,�I 1v�����!b���Wܶ�f$�В5=L���GmӘ6�+��`�K��x�^�!Ν��|����oS��ϧ��@:si���j�P�"tƅ�lW��Ô�*J`������PvM؈*�q3f_ �\@jd3$�?��fuϐ������jǁ�zx��y��9����ԼF2�@q3��$�/���9wkM�F攊�WV�����B�X���	Q�j����2��8b�d���7F�w�	.V�q� �#�:V�j����=f&�ʕ�� s��&��x�u�׹�l���S{�e�������%v��?�A�j�q�ʀ�C�M��k�2�F݌�
	c���9˥�����H�1���!R�<����I J�L35pm'�0nx��81�J��t�$ cBH����G�����(x:�-�z���i�I�'bq`�/i�*���$E fJS�g|#���uE����hK�d �'�4��ԁ�����Či � [ɠ�ф�(�F�r.>TR�;��
Y�wl����Չ�1���in��$ ٯkmLA� -��l� V�|�3��F{��2�K�-A�u�*�P#��7���7Seo��5n�g}�Qbj&��k�2,o�GɂH� ��
7�Ӓ�D�c%V��B�f��q}��H�� ��Q"ُ����t�
56�~Nti���xG&�v�
 ��m"�أ�4��t�̙#MC�/�ܑN$���