BZh91AY&SY�v�� _�Px���������`?6 c����M��&LSh�H�i���L###jO@* 4m@h =A�  `LM&L�LM2100���&L�20�&�db``9�14L�2da0M4����$D��zhiO�4��f��24i��C	��@h�o��H�	
�b$������@?��0`�"� 5?���ƈd0E��;�CH��ظ}��ԐL��ܖ| ����^Q�s�8}�+�ù���E �2��2��^*��^J--9�FƨHʙ��ㅎ0H̵i)���Z��4��D�/mr�K@���oQ��� 3�oJq��8hӤ?��h6[ll̚�w�:�uz�
���
�X2y��F�� �5-�+�o p	��.��YV|4qm�5$�h>K�^FLp�L\#@�� �v����H�H�d}A��̇yv�S#6��aPd�ep�Ĕ��T��*�CB3��UȪ���j�85��[�+T"Y��p��u�0�b����ض��=�Vʵ�MR��R���0�P&2��eTB��#��3�r�C֎���iFˇj��T�V���S��5��,ߟW��qA ��%��0@A�v�?�%/W��Ur�S�vK;nL�p�ё8�@�0B��kAAV{�D���b� 1y�*i��"��hat���E�F�*b��k�P�q	駣�4�+T����}�*�����������ND�����+�Fe�7�o��̦ȡ �4�(y6��uh��) ��U"�ʻ���JK��0@`X!������R(�d�=G fr��&��l���zP�SH�����9�\�ŝ�0�@l��7���;�<�����H���UT՞�F��b�y8�O�K
(�i��qZp�j�o�ޛf��!�/�_=���2XH\�
d��Z�&�AO\��dxi*4�Ԥ �Anmi��_��m�1���ұ)�fE��YQ|���_8t�":䎋r����
Q@`Hs*b��r�r�۸�Rݠ�.~,
I/��{a)�b�q�^IZ�>�a�H�6���d�א�8�y+�Y��Y�bnbt$��]�g�g^Gk��@�}@ꋨh<[
#
���i��3(��ŀ"���"(*`�8{!eR1
��*���eͮ���WV	�� M���(��$�2��sq�,�>��O�*p-���d�3E�n8�g�J��#Y�l�u�
1� ��u�i��]~0�z@��I���~:�.�Òj�R�9hVKf�r�~�vy#��8����େbks�X�Z��]TـXȱ�O�� b� ��h�.+4f�SrC�e�z0�6r��#	�	uH���D
�o�y}�[�gͪ̄�(*�Q2dp}�Ch�ʷf������#{M#������ܑN$9�9 