BZh91AY&SY��P	 �߀Px���������P��[�w�����ڄ�M&�<��M&h �D�4�4  ѐh4&�P��@&#   &���)����=OP   4$4�D��h�L��!��PɓM���&@OT�Q�S�4ѦCG�4�@@$	t�	"�H�J��'�{��$��~J���� j0�ം��XF6�V�(���Ϲ���l�ٳ2���;j�/���N�)bt#%v�%2�)S��#�oX����t��P���F9��ժ�F�US,�N���tr��HB1m!u���I���a����6n��R�~����»���؎=�R��ނ�ĥ;L��o\t*�e�;X�ɔ���惬i\х�[��s�v�*Pi��d��T��9�a�R�4n�3mJ�hP�g2/F�Ve0�Q�q��mL�ˉ+Me��)���!�Tդ8���h�R��j���l����^ݕ�R*�PuT�ob �,5��~��㺭���Cm����B���򔗟wm�-z�&L�v��Yf��\��v�A����(2��0��L�@��0���g�qh����X�l
�L���êTw��zq��p�K=�FE�Z���������Q@Jd84�	gC�$���%���WHf�4_aO}	��{6̐牌��5z��?)�e�9���0� �
A����vC`7ŴO#���ƵUJ~�IXY�!�B?�#z�Y4/��|h%����$���Վ'S$p�E�B�����$:k�5��ry<bY�N=1��Ŧ|���1\�Z�D<�ۜ�ݠҌ�X6
R#�	Ns�F6Af�(x#��ۑ1���AĦ��V��B�w�F2�z'M���Eb��I�����(�H��o���0)�\��H���Ő"=���IL�*���nb��1X{	��+|A��$��
1�?	�I�Z��;&y�� }S���v��K6�֬�TdbB�$���,�1�ZM�K��R=`�EV��S%�i�Ȋ�'BW�B�5.�jHE�e��'�Ȏ��7��×X�Y�TJ�$�N��( �S��h'�F�n��4�h�P��.�Q��N]~R�7H��T�*n�A峚��V��D��6hJ���@�ө�L��Z� yRA�{���o�%�����OJ�*��J8��J.��3�"�;�c�y\I����zJV7 %���Ĥ�;xFD���,� T�O)k!ƻ�QVB��aEZ�u�]�<�JD�BP$R/_K�W֍dKcb������Э6;������ F��t���˾z����$fi�]~v�UB���"�(HAӨ�