BZh91AY&SY��j" �_�Px����������P�8� �{��B*�$�4�<�MM�I3%4�<�OP�A��4~��S��@ 4 �   ���jz��2h �L��2  �0@E#�SѨ����L������"Bd#M(z��hd������ a1$�7\ .bD�$�����'�{W�_���6U�`����j��D�@`0E�m�CH�����m�Ն�	n�_��H��6�Km�x�r1i5TH�(\��٩�e��ԕ
�6����[$�b�	s>tg���(G)&��bc.��u�f�-IO5�I�^ٻ|��t� I�9��S�=���J/��Zv��X�Nɕ�>;���M'�>���)7ln����+0�C@]? �C3�Ѽ���@� Fڥ�%�4����[�D�dQbN�� �}#�D������a
P@i��@�.ͣ4�V��մ�.�%R�-��<�@�p�T�L���2�@�0�YQ�yOd��˒�.��(y}\	�1�B1�*�[�I|R�8xtD�Y!g"+��w,�C���;��e���$Z)�)r%`c����*Uw������px�UQE{
��A$��_v+�TG�ݦ�Zfr%&���Dt�+�J	�U(��B:��?d�z��p��Hֆ�f�}��xW����S�3� �،q�C������p�z�60ڃ��\�4np^�����K��12Y�\���%�f\��e6�!.n*��m0'��G���G����ʯ#��d{�s�KRӕ��;~��9w
A�!�_���\9	�;.Ŧ�A){�ρ.Vq8I�F{w�v_Ҁ�\��@��	|��h�t����'�6��!�W�~=�r�%('{k�w���W�vh%;igœ��p��v��	2Og�,1Gp	Nt��'�P\�#����(RINX�l�3+�����2���L�
I��L���j�#ڲ�[�_�B`a	=���z�BH�5�k��B#v�G������/��[
MD ��"l����։�6��	F�,35�m����#�G��4����u��F�%��[����`w��"a��`芐�k$*�EBz���Y��u%{ԽuȐ���RN�Ў�/�ӬEbJ�A+�I��W���*pq��Š��%���'A�w��P�
��z}ޒ�;�g��J�+.s�]�y�֤��#��8mJw��mt�u&���@6�	9G�Ϙ��O�t��2�+BX���c&��^$���I˴�O:_��
����<���*ʵ:�4c@Hy1��d	Y�J���l�Q2�A�s.Ye���_K`:R���A"j���^��nd0�=���ef$�)Ԝ����󀄫fGĽFv%��5���bɒ2��x��+���H�
�-D@