BZh91AY&SY���Z ߀Px����߰����`��w9 uqU�h)J��&�ѕO�S#j��i�i�OQ��i��&A�~F�ԩ @     hɉ�	���0 �`�0��E!@� h �  h�2b`b0#L1&L0H�!Oi��L)�=F�4� h=G��$����ڒ@U�I$$$=d%g�} @���T�f�(�a����ĄV6��*�����n|1�I�&p@\��MN��9;58'/VW�Пa*��2h�T�M�B bW*X�R�(���e+��d�^U.]
c��5B���\��V��ڤ��c�G
����2e'��5��e
�ܒ+V�0�½��ύɀ�l_��붚���h�&kfd�ח�=��/��4|�u�UFfIJ,����ޕ�P@�HP(����aEuq٩��M�r��i>�`V
�i���Ko���z�TZ3�ƍ�-�����Aiq`��M�#�ٮ�҃�(��b�Ä6d�Ȅ���8�� ��f�aE�8!L-��k�W�����RPW.y��uL��6��ا4�8�K�̿��Эʎ��p����")�-�A�[<Kn�7�ŕ����A!�@q�+��I(E�8`�:j+;w�&m_jtS�q�1h��KjU��V�b�u黔���6.�a�p[���+�af`ES��jG3c�3\��T��0�<T��>�H���I��̞�Y.NS�)z�m:\��ː�F�Ʉ*a.h%�Ҫ���³4x�a�����UEĖi�;RQ�]_�24
�q���30$��W5���f�f�+q��G'�sY3Y����X:AL��ghm��k[C�����a��^���6��{?|~u�� ��IEg��u�j��=���N�Y��Y�ge�J�@�^�f'�5�	qqD��/�mP�{��! ��¦X<ݱ����������@I�16��ݱ�qk�����͋U&��o����K��ߝ]����*Ld����zj�Du��
�B��誃v"��v�xБ'�K��:~�3P >��߿?�y\�`�!}��946̄�^��=��>�ǍJ����r�X��qG��Q����}l��.� ������G3���D3	�\�Z���{�X�����%�Κ^����v��1{�t8���{.p��Mt�(z���A��4�K�d��A�u�yJ*5 Y
��L�yn�2� �c+��4I7���������4w���)��u��L��,H9��F��Uװ&>�b}����\�N��^����?qSp�_0p�,V�k�L�8���0�Z���e��ճL+�Kr�1���h�sI7����]��T#c1��|������H���jcEdFbiԕ�Aj_bHD�e���g���5gR������3S��* @B�G{z���;K ���)�NT-�Q�{�g�vD�-s��z0��dd����i;��b�l` ̜AI�p.\C@=� !S�����[f\�{�Ζ@�c�*�P#�OD�5����-�p�����*c�ʢC����ʏE�bEN���v{\���z�TFfB��1ʬٲ]xh�~���$9BF)���<��}J-[�g �]���UNFm���@b�>G:��w�V�6{"6��0��~<A/���)���