BZh91AY&SY�f�� �_�Px����߰����P�9Z�G8�fLf�	$& I��m51L������Sj���P �@2 @L�DM5LFM4dچ�@4hh h2`LM&L�LM2100	Bf�L�� ~��LO)�d ��14������J�$P$�@+ �	F��P�����P��R�&��밢 [�HcT�ѵ�4��Vח�M�Z���%��@w]���y�٘�Z���n"fB]�v����TCdٶ�8L�uSӹ�����:Z���*��8�p�8$3=��'%v�ͨ6�pJ����^�Æ�|�>��B`����V8���8(7Ͷ�t����o&X�7�'�l�컍j�R�����Z�ڪ��ӑ��x���Ql�^d-7l�m�����ճ������:	5�W�[A��r��β�9F���1'WZX�w6Hm�$tI��.@j�C�l��0rqP`�e �D��UAE� �^�e��4EE�I�w�g�Q3�p��k.�\�f$�����
��/�F�6M�3�^fJ$ĕ�d�Zi�-�^oZ���n�OY��~��m�M�w���K����-Sވ�%���1���V`ȴD���1��(T>��mP�h��Bb��7:k�X�2a[T�,�%��b�����Ȝ������������A_���>z��_<�H������r,�4!z]��ϙUْBb���L��Q�w��Ƣ����{������cX�����W��|ۨ>�-��8�B�7��Nӕ�8����BT�	��˸�=�B7p��_A�Y <I�B���c�k'E�tt���_ZC=�E+���JpN�R{�'�[�"�C< �NCs�e1�!�Ő�A�ĦH��N�94�Ⴀt������!	�9W�,3s��eSݪ$���T�U*��B�������l�r��}O $(�8*�+F��QՈ@n:HwL��ɂ���Rj�4ы[@t��+�paN��B9��lc�O�H=��+7rS:��,b���8 <hB�̶|#S5��x�B,��#��oh�2�D�F�щ#d�w'6 S���",(�Jp�pRFb�Y<DR�M�!�D�m�y��Br�A��ڸXfFBԄ,��H=��
�^�����a�3���%B�9ͯ7~�8*Y#I�5���]hB~�2L��e��NTq��y{�eGn��T�J�뚶��P�;,4@� �呌0���`��~pR��IX��.�I]Fi����Ski��d!F��M��r.a��Z4���t�m4�ڇNc�@9�$G�����Z�z��9T������ST��6�py�HV���5�$�����u��Hœ$ci0	��ܑN$#Y�(�