BZh91AY&SY�&  _�Px����߰����`?M��@ABI"O�b�����=L�� 4��S�T�      4d���`F�b0L�`��F�4CA�� @  4d���`F�b0L�`��h!�z2L���i�14��G��J��� �(���$"����G��_`@y}�6Te�TC���R<h F#Y����4�����%��N9�40X�^�+c��+x�j��d��ؖ͠hD��s0�DM��d�&�46������-�u��2�Y1����$f<2)&���ރ0Y˔���D	b/�ǩ��i�	� �{��]}�ʫ��ib{�j�y:(�C��.�\1�M�yÁJ�Cx�}X�l�xKEN��H �PK ��o[B�ɖ����"�G�'#���Z��1�r�;5#���L�����
�pe����Yw�c�{��mjm��S
8��n�����,��1�8�i�$dɃ�0f2ԓ:e!	�d���!,g�Z���0�.U5$���;���7�-��k��٬ݧ�5��#z��X򋱋6D�`�D7�ϑp�DVw��}6F]H�}Ά��r�[���U����}��� @b "�m{T󒗳��Uu+=Qd��Z��K�^4���h b1c&�]�0j���!eH�@1v�������ara{U�(b�@�0��J��Gs����$�[��3.�:$�6s�&����yh��#��|$���k�Ҡ�����1ѨHc�9�o���߯�RH��3J���p�|o3�JKW��?���}�]��:����'���|��^�U,=�$�p�zN#ȋ��uv���� 9�f��œ��ڈډ"����6X����\��o�����:���W������Z�?�ݵ�g�H0��b��L���N��LԂ�XqGQ�בR�"A �1n])�0.����l}��SzLKc����{��]^��̍��B9�~���2�.$9U/F�lV��
�YN��Rט�.cg踽eNa�ް��9-7l�](
��cc�{�� >�8z�����ݙh���0�!����v.�4B9�q��s�b>�uE�4IE�T'KlcE����7� ]gd��p�H� ˌT� �|#}R3
�Es���h��&�%����,!
��u䘥AX 1�A�n�8��9v��/�%heu*$�9�]b�"��0�FSpɎv(����u&K�H��C��@B�M��Ȼn|N�^��%�;/Y�ʁo��R����m5V���Ͷ��}�侮3Z䬼��U�q%��g{.�9Z���VS�K�3������5l��E���(�l�U )���e1гH�A��{Π��PYc�<h@gm�V�_���-�����4��ݨ1��ܑN$x�ɀ