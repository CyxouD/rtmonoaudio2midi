BZh91AY&SYS�� �_�Px����߰����P�ꛀ�8Ն65BIh&�)�I�F��26�F���5O�LEH�  Q�   � �53$ѵ=OC !�j0F� 0`��`ѐ��&��DI��G�4���mM?T�I��h#A�L��#.��$U�I BBWH	?�������Q��6�C���;�$,��G6�*��vo\;zr�q�넖w_�
��C���:���=>x\iΡ�BF^�C�8�#�fl%c���Nh3	x�HB�9H�����8W��{�7L6�ӧN�Ӂ|��>��_Z�:�w'fh��E��pwInv]@Ε�ĉ�A������2��_�h`�J��5�{kq��;-�Bs��fB��������3T����h�v�:�DY�R�a�f��`�� :�$��"v�Pj.��i2��3T(��5�;����	�C�zf�écSy{,7�Z�=K�}[�K0�B��-,��k�O����nRH,m�m��4�	�䧌�����Z�g$E��e���M\b��!6�ٖ��T~ƈ`e�39��!��px����.�i�7��l���޽��^߁{e�=�ٴ�\S�{q�	i���������;��,<��ё�2��ޤ:�����)��b�G���7\�x����<h�T��?"'�{^��ʭܰr��v�A��)�C`#Ą����n<����T�gVM
`r��p��>>��!��<e�'�K���c@�j,F̤W`R�gӛ�Z�m~�8�N1+tQ�zզq��4���۽3�P�^T՝����+��L�L��xay2��G��K�6#����*a$9̯{v���_����A�1�Ϟ)�L�努��� F&��\&G�����C޵'���F�M6u6{�p�!�$��THl��&RV�"obl����c�>H�h Dj��0�d{`yz��"9�r�2�b�+Q����!|�G�*��#�t��9�P.�:��Q"�	ն1��F��7hB�5>{hH� �*;�uH�����0V�PE�D���yJ� �K{|Y���g�	�m���CU�!���A�#_;����3X�����6��#��}��╥�?;�F������&�`� �)���9�|	]��N�Q�eJ��IC 3A'�5D"� ��th4C$h�I��2�t�O-QC�M5��8�}!!��z@E��=)���X#�����WE�J��E�å!�:Nd&�k�%�[���?,� ��++�6����wQ3m�j��K�۞�ls�.d���-�B����)���t�