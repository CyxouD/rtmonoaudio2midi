BZh91AY&SY��i^ �_�Px����߰����`������ �<�AE �A2�
4��4zF���42d�5= %*0       2d�!�@2 Ѡѐ � Ф��       j��@4 �M     DD�4dS=4�z���G���4�2h������ 	?0~ay���_@�^����X&����(�a�AX�sG{i0��\W?�^:�W%��]='��^`��|�A�)@��VI�ѐ��2�) ��@q�) F4���%CL9�C�� ö���i��q�p��	�F��je��T}�4
�9I.�� �^X�e��i����lo��j��djo�y6��P|4�5�b��Ў��Wʁ�\Q���%cH!))^D*��+K�U	m�����QKE�Xߌ�	��&���Vs\	m6��ʲ�l����* *R�2�jPx<<%B)p����wGxD�	4���Pu�S��M3c-S��J�pB��(��D6oJ�*� :�p��6�P)UC#� ��P��G��p*G��.�`9qa]���"!aj��hK�^C�@��I�I0���!I�2֢��2��iP�=�*�R�p�V�F�.���`9{!�]�`WXwI�b͇��q
 8(��p!�b[v�e�ٚ��C�Tm��M������ �b[nt�Y��U{���i�w���^lH��h�2�����U.�u8�뼯��N�=�W�yJH � p  A���b��'.�sG��P�@	�b/`�m���0�%�ld��4*����"��1{^g��[HX��a{Q�11���� �[6/���/�9UW�6<��J�����B���w�)黏o	�3	gҼO=r,�өL.5���eX1!b���L
;(#�f^��-��ZZ�}�B��31r,�$����C�r�D�c!�.����>kS~��,�Q��'<~G,�\��:2÷F��ϩ��X R�K{l��Q�M@Y�̱��CF��nÄjJܲ���Y��i��ݟ;��~�wWc?@����I
 �-)�+��R
p��u��,ʕ����u�j��q�y �c.�����TQU*���
�8��(��`;�rٙ02'�89G��	�m���1����Y0\�������D�1ke��}��b�8k�cc4����¤N>���7�@`mi^�@�}k�P�����s�b> ��k%ʪ�5�1��F��84P&��DPT�Jp����`+��UM����nQ,��K� P��������dl8 Z�D�s_��(_
��<���1M���oS�Ԡ�����x�r]#i���ZV�0@��~l{���\{X>�@�W�t�{���9�}��֖A���*�P#~��*@oC�)�c;��^��p��+ب[!=3	.7��`@�`�]��*��UQ������V���9�a��"����Eُ��ɋ䜶z�ĺ�g �ۊ-RSr3a.��� V3#�fQ��ǡ�ǥ�H�ɒ5X;v ��.�p�!}|Ҽ