BZh91AY&SY۞�~ �߀Px����߰����`~��s� �}z�PD($���2&ȓ�Lh���2mO(�h��!4�%P @    T���zL&�F�dhhɦ�� ��B�ڧ� �   M4j�h��@    $HF������Q�S�ʞ���6�2���!	���B��` ��"���=�� �O����,��E �0�d�@y�I#�*��Ʉ4�����e�� ����P,�-rZKFw�M�n!�ut+�  @5�HR�
NPw u5��5!�'v�3��o�Î1��4�!M[h��;Yc�L���dce���� ��� Aj�!$��r�5Q��<.�`3G����x��/>��kZl�Aq��k��ͪe�T3E�܌�0�Oq��`TJ$1�^l�G�K��l�c1R-i͊/��
�@��7�M��8��-��V�-�_"�Eed��]S��j��e���s/Ĕ��r��D%	zW+�EB�weP�-���иu�������HS0)0���t�ת�D���G{f%���k�)�T�u��_U%n��3).��2dh������	��Ob�b���K:�����]�m�RC�<5�i�e��,\�F��Sp�N�Kov]&hF4L
��j9�(�NU�IRd��,$�����݋��f�����`��	W��Kr$����Ebu	�t�Y�g��m��
�l�@�1���BDE@�ɅMrsv�C&5O��1�f���r������Ɔ�����DC_�@;ǻ��^�L�ӑ�Ma�\ �-=|�?�!�`KM�+�R�7�m	���J�)���N�P�c����8M�}CȂ�E����<�@�/O=s�n��E��Q]o7P����ڗ�c͡��`%ڗ{�&OB-�E�qAn��FAY&��3�"S�}�JP��T�v�L�l�`��߉o�[�q�3
L��b �#���:_#�>�*�#���td��]��2��y��A�c+��$��`W�T����ϐo�DvȎ�Wv���)(�;����u�	��A>3%��`�W��e�h��e�8��m�
�4���#` �c���<��ϟ@>4"W�v���v+(�r��C:��ܽ�e�gm�s�"a���!��̚.��,�c-"2&�I^В ^Ä�?+�$"`2�
I�3��D�Er���)ZSPD�	UD���xuxWT�6}�# 3�#N�H7�Y�Q�n�=~3�8L���PAK67v͏^��6�# ��l6��X`6jnlLA��-�°m��_�����-�N���f�!��PU��F�~�t�7���6�:]���A��+�I]Z�V^��pT����/����"�e2t�`�M0��*\A��Ujբ�Ûe�?Q\H,��R(�lՁ�Wl"Yk�:=8�	bSW�3:��<��F��{͊�e�}�l�H��Hݠ�9����)����