BZh91AY&SY�l1� �_�Px����߰����`\�[��5:4e�A$�D��T�T�ڞ��iL��&ODz�4d�5O�R� �� �   "��6MC&����hɉ�dM�		����i�=OP�d�M� 9�14L�2da0M4����$PL���L
z�MI�<��Th@�JB��y$#$Y$�Q I	I󜫨ߞ
�Ń`��5~q- ��$�p�1�y0�H��Z�q�U؀#U-Z�
g�,�_m冷O��
����$�ڇFln�J�j���N�9���8Pǉ�����	������ ��Ki�m���& C00x���m?����n&�eRy�;p1�s�xu@d��Rr�ijI*i�)��j�kK0��mL���)��J��10�et�TE��q;0.d9��]Y�Y*��;�՚c5 Ӛw��B�N��Z��$X"��T&���)[I�Jb�iZV�0�D3�����\��,2�T��!�!�)ˣ�lW�Zef[g��ą�L��Jʼ�ʇ"d�}���0�/������7b��DZ�J��r� ��X��Κ%�S�t�hi����$:X+����[l�XCY�`��I�UȸgܔpH;�]�Jk}
k�6�`]#����{����~��m�@"�8w�w
K���u��Z����	/s����Hhr�"� cG0�4��6"�sM� ip������0V��­O�f�4��^�e�xz��A��uDO�Z�>3 ���b������Yg��@6S����)�* ��^]��5ڀD�"�B��M�1.y9�$Z
$X�q�wq���z�0�hm�k�+�U-�#��`7�A<ow
��=(|T�<}�Uq�#�t�+�N+�1�����ʗ�φ�G3&�Do�D��+�ѕ�"ֺ����h%Y(s�m+�ǥ5�\���g�[,��#F� �'�
��X�J�@��G�i�`L�D7�k�3+Jx�.�d1���"��\Yu��!>`���p�-��H�:wq���@"RPdV�+Q�k���=#� ��a_I8.;����Ws���d���DpZ�ݜ�6 ��llc�/�����ۧI�_Fq�e ��I� �<W�A����8���4P�A���%":��х�Y<
ɡ$Ay-+�h�"�35I�g,Gz��Y<d��R��B�R���,��C�/���ޘ��� F�eB�ZV'��5�|�p�9�{7:�K�RX�5������H� ��ÎLU���!�p��f` ����{t)��]�'rԕ�Ϋ��M(�Ձ)�7� �>���uN�Xa���t�+�b����\S�;B�K��� EX'~�A�]�qL2dT�@�r,Ye}m��s�!Z�
% �I"�ݚ_��ȑ�,��rs�Ej
w#M�8>o@"�d}*]C�v������ɒ1������"�(HJ���