BZh91AY&SYG���  ߀Px����߰����`�' F�R5�PI �	�ڞ�
����M4OM50�@j��e)   @ ��0L@0	�h�h`ba)�)�&��h�� i�z�    �@9�#� �&���0F&$SU?I�#�?Q�H'�L�@4ORʩ�� p��E@�Q�hY�?g�"�/����1� '`�F�`{�z���s &�8@��2�O;��^|BD�:���$�N[z��XYݝFrr�2aUPAD�TR1U2�1e�!y�WM35w?͒qkT��1�Bi���g�S�tX����t�uL5�CP^k�EC0�`��|8z���&���w�=�z����8[�tz<M�y����9��=m�A�o��72���ްTȃ ��Pt���Wd�1O/�i�)�4��Vlm� w8H\��6Cs�V�5)Hh��k�"���h��eu3��gq^mR	�c��z�'l�h�Ӑ�"��6�X�i���ڹ���j5��P��z��&	��a���XTj���B�+T^Q�*bdA�;:�)�ٚx��-�
���FE�t�@6*j�6��c�P)D��.��Y��d5�5U�4� "�XiFK���\�)rl��˦ehi����:���4'�|a��U�6@���J�}����,51��#r��Ի<���!YCާ�-<Jz�X��׃\M�^�?'�ܨ���UA�"	$�w�q^R�<��n3��l���f�8؃R�t�I�Bd���G�4@��$Jrfs R/�N�8^�x��$���6�! ��G�����a9Yg�,o���^���z��)��~��W���쨼�mzt`[�b�����?���,���,����U�Q;��q4hQ�m��3�#�s��!#J�㫨:���v��#�sD�E>u S��i�����.LRUv*��W�8Mqі,�/�]���B%ܗɎkF�s'T��H�bz���r�5���w_�JpN�R{�g���i?L!NI���!�z ����2"�TtZ-�-�� ��T�V}-"E�!!�B��L_Y.%���1*v��L�YZ�A}zD$i4yv����r�M�l���A�R�+l�uY*�� 7F�3OKU	��O1a��=DNa��Po���%���r�#M,36���Ð�%[O�~�����N��8�=�����t�s�3�7KR\3'8M	�Q���-��"ab����EA������CA�fP'�`�q�j���f�9�&��$�D�s��`(�:�yqro�lN�r��b����aM���w��5f�C�����9��:�K�S���ξe�Ђ)c+m����a��x�A�6b���(H������wFš*��`�Iö�������Xh�{��[�w�R�芲��ڤ��z�	�*6�sT!"l!"4��I��E���.J��:�FU�9J�"���s�SD�ؽ�������`~y�Cm�ʮRSr2�׭��BE���2Q��c�ُ���&H�k��b���"�(H#��s 