BZh91AY&SYj!k -_�Px����߰����P�b��%$�F���02A'�ީ➉�=F&#i���� �� i� d   0`��`ѐ��&��0`��`ѐ��&��DA&�S�d���b4� h �)1��BAf$Q %0@"���/ؐ��ʌ��b@5>�e?#�,����E�`���٧����޹,��GM��o(vk\r.N8��R($/������)IRPf�2Ɏ:�,٠�������E�A�P -\�Kl�9���>��L$00y���N�'�J�4��QS���܀��'X貺��o'a����F��"�ZV�A���QF�d2ӄ��B��镂$p�̪v�V�la�m�@�`��|����V��%�ō��&&S?�#��Be�*6�*`�;6l.V��4l�$!8ҡv�K}N�9
�  �WaR&f\�E:V"��-�%HhK4�% ��{K8t���T!��;b�ć�I{��u��yJ3Uh��#Zcy$Y��Y��Z� �bK�47L�BҸ�h߭���JFU�F��#Wn�p�h�D��P�Ɋ�����|���	�1$�@:ր�	�?mO����8��J�E�,��ׂ�3��Z��+A���)�l)���H��.�YA�H���.0����L�d$��X�Ƶ��;�*{�S]}y�Ϡ�\)��d�	j�g�����Z~??	��U^�vBފ�)	�<_B��IS��<��yPG~߿�u���`�ρ����O|Am$im���20~���Ep�hlH���fr��&���n\�D�z��!���|��:4ϟF��1�Z�.a )�KsMwl�J6=":����v%fOr�%��g;��JPN鶚^���7�&���Z�;sSS:� �(b��h	��ZR:�	1���%��:9O���UiH�r-��3Nb��amyv���Jf�VQ]J��v	Q��`�ltӣnt�� ��ኂԣR(�B�F�����zY�$�|�
�� ��"l��C��d�=�6fa�a�{bzrvDs������x2��£���k���܎F9�7��"X�A��Hh5+�P�M���4N���@��U�"�2�
S�gT#�T���Q;�U^%A&�%��u�XI
���=�,�єH�@l���6e&(a1�~}��Xdm�velZ^�6��l`�Rd�A��:�fb@=��Ў$�p.��P=� ![�y���)�ue��G�ŕ+C�R�oa����r\B �"l���f�X�`�T�=�T������t���,��-a!�5M�L$m�K4Y�V�����G�9�*�.��mC�!�JN�(�m7��\��м;�g Ǆ���IT�h�׭��A$���n�ݘ|��峒!#}����9�?�w$S�	�"�