BZh91AY&SY�G�� �_�Px����߰����`��,��q����AI&��)�ͩ�L�z&�)��4�dƠ�?M �(�`	� `	��ш1�101��&$BS�A�����h M�101��&$PL����M4i���O)���@�	�DXH�I 8) sģ��/��#��a�`��ju�p/�I �"�6��i0�^-��͢�P�w�;����v����Q��	��޶�j��|%����cci��3$K-U.mgV�RLL��w���ӝ�7�Fe}0�����r�y��k!�r.� $M� R-����<��2�``��֜x���j�3?͉40 ���kƽ�ɮl�,g�Z����F����ͬ��엵\r�����mq�x�GG���z�n�Dr,��C�]�%���y�Tp�����2�$87��d=J�`��|�K1�D�Q<��هzd&����f�]�!�J��u
�̂���M�Ϲ�2Bx
��N�S�܇'�3FmroW1Q��ְ�vפϲ��Y.�)��,� ��U;�>�P�h�Ne*�Y��̒2Keda��L�jYv��ؕ�Մ��w&���i��nE��0����P{�
�}g�����X�f�zSp�gr�6��øM
�MAs���}ޟ���BH$|��$"&�^�RR���e�e��lT��;��/�����Rn �P4q�4�p|�%,H���EЄ1r0����4���Z����vCa{/fO����.���z��5-2;;�|�wo�xyn|��߷E3�J����,��q)!�᾿_� $!�i]�|��p4**z�Ns��Ni��c�od�Pj���r�D�3!�! n��'�����ڸ7Qt�̢I���Vi9������f^��@u�h�!�ԼX�ńs45
#�)�(�8�z�Ŭ�5�C��%Y(ז13�e��ӳ��j�B���9j����ą��F$:��4�:ľP%���r:�M�Sj(Bo,�$̭)��yPb1��Ӿ�k
H�B��y�!����##ǞNi��֘1!��uA�9Tj��f��`H|5��E-w��V��>A���^B�h�^���V�poBÄB
�a�a�{^{o�t@s���
e���pL��u`l`�nB��\�$������Ph���D���CLh���Rw'3
���I"(X̥8{aVH�,ʖYN&�rL�u�O�\0���|�,(Ԅ#4!<J �ߨ�Sq�Vx�W��R3lv$��͎�k�`�X�#� ���ܕ"Ƅ!�x#�2.���B�����+����grҕ�«@M��!��q)�$�y�ih�wU�����wLMZ^Bs�X��M�P�a�^tBkBf�d3�M2
4 b9,�������H� pq�$G �6��`Y���vR�A}w�N��pX]s��a!���p�Ɋ?x�{1��$\ɒ/�v�LAW�]��BCm�@