BZh91AY&SY�� _�Px����߰����P��4衎��VZ�P�D�&A5=<�)���M���@i2z��Oi       BA52�z �L�����i�4z� S�4d���`F�b0L�`�"
��~T���5Oh��@�h�$�,��@*X�4$!%Z�HJ;�ù���~XT̰l�j0�;�H/e�J��)ch�a"��ϩm�b���K
���Bݺ	o�u:��-B�]��*x#�N�q�a��0�|0���9[5b�o�#�qkP�����Tj���|�7
t�	
W��$L]�j�=�<�C00j�~g�^�B�Κ�3g~tz`y;4���5z�%�%���s�lݻ��M�T�J��v5#QG͸��X���4��Ƙ�č�%9�Y@�$�H`e����=c�r2��6��Xy��pr����զt�i��C3k��ʘ+��:o�0�<_��1���7l�)oRCK2!Bi�	F�������y"9�}	�Fh�޵�Y5i��ګj�ݽ�>��m���Sm���"�|�
�����]7Y����u�{��i�kft�D1�[4P���
n���"��as�z�y���)��_�\�!�j1kf�w|��J3���{����'w��Z�~ߏ����x�yN%�>S�����HB>7�]����a�19��ʊ�U��ϧ��:(��~����"�c�!=Wq5>��B�EasCb�B�y�	�=�����V�;��?C���G��r�ѫ�~�2����`�K�/팵�4:(�������P�X�w�g;��JU'n�1{�V�E�+Z�D<|v�gm�Ҍ#��<m
��p(w��oh[�~H�4tp\�B�B�oL_a��W>�zf��\�U����_�lҍr$~!�N�d��"RP��3����� �m�J�����>��A�Y��C.g0a�d�Z�U��|pB(�#��~�q���պ�9��pXid	k��������υ�C��0�{�Њ�h1�ESS%�cF(��d�V�$(&���1B,.�T�vļ�HжVYr�V)�T�)&eu.%"B!P�U@��{KьB3Fނ(?����Vʩ� ��~�@둳�܉�(fs�,ގa��4��#�o<[R�Lb�Y�oL�퐷m�ڄ!˦<#TN�2Z��Ǘ�YҠp��(c&�\	�0n�i�x��
�w�Wi�@VZ�[j��G��-����X�]�U��f���r|GQZ��J��f1i�(�H�T�i�<���Z��L�;�]�l�I]�*NF8�8<*HE����E�x�����9#CM#]�t��ܑN$iG-�