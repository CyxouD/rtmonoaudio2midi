BZh91AY&SYHe� �߀Px���������P�ޓ�cx�l�JHCA4�ji�$��FSLLL��h�h5O��@с4���#!���L�"h�Ҍj4mF�=&��h �j��   A�  "�zd�#�Q�=F��m!�@�h�=t ���I�A?2��i����L��C��6W愅`�1�s��H�
5��p�g���+^����n��u�X(伭l�	��7Q0uX�7?M�UJ��j��c��YA#43I��qm�3�9�\tqHB�*�$"�o�6U��;y(�lj�~��.�w�q:W��X܃{������y^�?�Q1���d�%��b]"���nr�*�VF8� ��"e��@@��t��;�f�5A��Q)[P�y�k6�F����V�6_M��X�T[�J�
X�M�i���"Z=(�ԼU�E���R3/��
�F
T8�E��2÷X��؁��E��QA.���Hfe��������bX�����lA���S�J^�/r��i��%���x���,D��a��`���0����� �.v3�����U��aF��1f���kV��=p��JN�7[�����c������S���|v�����SW�6<�1V��Q�����(��b����q��� ����T�߅]d��*�9Ɣγs��� o�{^�L9Z�7����m��{:$�}I��ʽ�ّ�$��tp/Q���"=�"o�1Ø���`�r�nJ���E1ZՊ��qXҎL�y��x�4�U޷楨C�ߞ���T(d1b4��L�rҐi��I�\��R\V����y!�4�n*�����0]"/Ѻ�=3c(%�u*����Y��F߀�6�@��`�DB�tK-�[t��ClA�g��-�4���'1!�cgW@}K��%f�$�+�c���06�>~]rQ�_J�o	����Ĺ ���Ǻ�c^�r ��r�QzTN�lcFF����Z�MOM��"�e�T� �l#]�2*��YM�!�Y��FB�Gk�pMn���Z.�� �!X�|)�@�r�F�������),s�E�׌�²�Fa��5��V�C�݀�Tȸ����@"
~:F���yaa�G�\	Zh��1�5qh3H!��:�-��F��S�5�SF�9H���j��'	�*8��������C���� �2��T���V+��B�"�̑U��=�K��@�M�rW���;��a�K����u���}8tųl �������?��H�
	�w�