BZh91AY&SY��� ߀Px����߰����`?z���s�0P*�H�I��&i�i��mG�d���=M��j����P h�0  b` 挘� ���F	� ��(�� SOP�4Ѡ z��C�2b`b0#L1&L0H��!�ѓMM�S��M6� 4$H~;@As( B�B/��"Q�x�/� 3e�B(@�1& :O�L�*$�b0E�m!�\����/O�V9��j��!N8`Sn:�U\��N���X���)��L�䖘P!�;&�	�0_r��D_M1.ʚP���z�!Ra4�1�f�o"��u�JIy`�x{� � Ɂ���z1�5t(��py;KR�]�.�OW���g�3u�q"���g"|m�Gu[��N0�8��� NĈ&�T����c��gw�Pt�h�\+we��@Ww�xJ,���,!c<S��)�J�&֎����+`w��Y�j.gfNB;�{�Вj\[�87�œ�)] F�b�L4vt�m�n0�M�Ӂo*5Q�8��u���TL'"2�e�$�4�5	 0��P���^�
�D�{o9���Ȧ܆�p�uY�ӂ%�1�֞B�ĥ��~qc5BBK"I$� �,;M$3ud�v�i�}�H�V�<�Z��3��wu�"`�i*3�b!�m,YVeH� �0������&�_�k|���fN����>�޽�n
󛖩Ϗ�����	O�������_
`XU�M��g99�Ƞ������yU�D �4���	�����G�:j���WU�t���Ac1�@���*P�;s1p0&`��v��<�^��kXlD�K�9��W�;'G��gDn]��:��܀x�����iK:}��4�s	�Uv>��-u^��G�bW�G�i�W�3ﶧi�U���)��
@��Ca��CIL��ҐiָI��S��(�`u�T�� 9�]�Jf�z�+؃1��])�F%�h�YU|� ����Q�$��;]�b`�2�;��kSg��5�	ӈ�� ��R@^���H�l%:�f�C����[f��:� WG;���� �T��Ǎq��7hMia���րR�@��}؞���"���A�!��J-j���4ƋI�N��Đ@��;fH� ʗ�N�p�ʤ`+��UM���&B	�D���x� �P�ٯ�=�s*�d l@^�ts`+���<�����!����OAI}�h��nJ�i#��{w�ic@�c��1��s���.���$��R��m��W���=X�`�@ ��;�T"(���j����F��<�~��A5�J���$�ߖoe��@�gJ��f*���Sb�B�N��{0��}䅀��Q"�լ��;x�9�{�p�v{K�VW�6j6��P@6���V̿��َ�9",�#-C����w$S�		M�p