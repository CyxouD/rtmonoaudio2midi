BZh91AY&SY/��� B_�Px����߰����P�s��AǮ7:w\ܬI	�SȏM2�bOH�<�mFFM�E< �� �     "	�)�e14L���   %���4�C��4 �@h i� H�4��5M=����C'�z� 4 A<�qF�S T( �t���m�����@�ʤi�s
Pz0Et�Б<0)����{<��u��*���8��<���ݪA�P�sI5�61��?�s�F�T$eM:X���cH�B�4-���ѽNn"��BH�^;�>-�é�Hf;���-+V���k��<�q������tLCTJD��^	�"nYPX�M�M��m�r��m��e1��hl�扌�$X�<�^f��Mk���E+��X�Y���ZH�e�A�IwUgG�Jc���B��d�%X�9P�Uh�D�X��:D���I��@y#�)WRTPg�Wo�bT�F���,(Ec�j�R�Ɉ������ ql�`Rb9FI'y0��5/���>P�" ,m��m�A�_
��J^m�W)`�;�d�����%�fa�bA���aTp{�K����������<��aa���گ��60�코x{!�;<����B�ص�v�sY��G�QxM���~"]i���&̞�G
����'�h��By	xJb���쐈i))�_>�y���b��Y���s���/Z&�*�J!%�(Α�6q�٦�3j�a�G��ޏ�Ks��Ŵ�<��I#�����T�SQdp�Ew�+��NeA�0���FݢYQF������y���M餵K�Wu��@Јp�����H4�\I��S��dr�>�H�ƪ����m��/�3z��fB��ƕ[�\J�T�K��$�J��o*!���=i� Q��XD1UM�Z���]֤>�Ip�"�:	����y98�̘��b/����ER�[l���$�]���Ǆ^g��d#oz�g����'=��[RH�t-�rA3F���q�*�����E�UI�4Ƌ���8`�A�}�̨�L���z'*h����J�(M�K5;�`B�GM�>�]%h�$�RHϬ�̶}QѢ@�������?���H(f��l��0�R��#q����b*��W'm�e��7Bp*�q�ly�E�ƭ�����V���Vgɠ���@ޓ��2�
��_��z�VO:�ե�')QX�Z��й�cf�s~ꦈ�[Y\���3�ܡ�uZt�;Cm��!9� �n*H�� ?ʕ�A�:�l��m�bX'���k3fpo�T3#�j�Vݎ虍NrE̙#
]����.�p� _Y'�