BZh91AY&SY(
߆ L_�Px����߰����P9�.�F�X�v`�A��i��4L��6�C4A��2i���j@h4  @  		H������4�4 h��& �4d40	�10�Dh�������i2@�G�� h�!-?�Idċ$�D�f�I�%����d��0l�j0�ം䰐i"LmXA�I��s�.^ݘ�*�6g\v���y��u�Ε�W���ؔ�����J�Zu��ڱC.j��9�Z4B�=$6��'Z�\���c�BD�|D��]72����V�l~�z���n����}�ף0.��=d;�-�ག\~{p���U���6�2��P5���p��|	ɠ�������6�$� �����eF�N("5�'&T8���B20�uZC6X�����i��3D誰JBЂ�q��J��x^�M�|�����D�7�m��4
����^�R^����2��L2����,�\犫E����j�P�-RdiyXd�C�hc��3j��20���,T�v;�S�%=s]��[z�˫�����*��y���7ۇl�f�}(��8��ѡH�O��Ev XP��&/'�LG�J^��y���V�8ʁg]��L"�~�� �`jhl��`6r��&����+kD��3�B�/Q�tx���ud�^C^��X
~ĺ��̈́h��t���'�V��P�]%��g;��JPN�T��R�÷)�k�MD<�V��}� n4���$HoSJ�����x���pi�F����E��L���^�|�<�~(1�d�\"�����RU.��)��:�Hs˽�`�(�b�QR�W4JW)��(DnW��z\t�����HAc�"^1���Nx�b��#Y�F�Xfk�. nx�|���w3NEU"8�H4 ��V�)wY����N�,G���{;���i��k,�EhhA�{����3T�|";7H�,Ֆ�ĥ	`�d�3m�p�A�9��=5# >�tr�+4B�H����*C�#OS�OAK5�se�ݠfj�H���Æ4b��0�'2�2.�:>`��	�}�|���k��v�б�Hk��@�1�;?�(@�{��d+� .�{I/׌��<��+V���$e$c;܀V�y���W�����è��2[0τ�|�-��X�QRD��5�y���A�X��g Ӻ���RX������fGq�Fv%���f69��2F������.�p� P�