BZh91AY&SY�*@ _�Px����߰����P�97Y���U�Ѣ5=)�$�EL�'�2 ѐj���M  i�  "��L������2� i���0L@0	�h�h`ba"���d�M�Oi�M�=&�4 �4�i��Av$P	
�d$��9ʿi t~7T�0l� ��6
�=X0E,m� �)aS[�\>}Z������,��N�7Ku�WP��J�	�$��n��s�#m�$fWթ�5�Zi�{���?),O�� �3�$ Ћ�	H]4���;�I� �`�y}�ٳ���[���9�� ��CY�˩��/ dK�.�z��-&U-͹B�M⍴]��Ĩ%X)�DF�L��������ib^��6i���2�d1S5<�3�Jb2֩oM-fY��l�l<�X�j�ǈ�b�c-\�L��]�Q@�C2��9EL@������\ m����J�iT��,.b�ղ�wG�Q�C���f���Bk��5���2�Xh\[��Y�l5��P��	�ª ƛK��l5���q�0�B"�B�	4��������,��|�u������trk������6�l  �oú����|^+,U�~"�pDZ���!��0�@�D�U,�NO�
	��hыb�� 4��R���킭��5.p�$�
L��mok��F�4UW._������n�}=�%��y��O�ۺsٮ��\6�Yf��T��n��,yK��<�L	��&ݫ��a�M"OXU�{�o�K���Դ�ot��C���A���@�lܶoVq�~5v$A(���9rt#�:٪��f�?��_R@u��϶7F��4m�D�
+oV7�H{��_��o�%'k���Uq��f8���Z�n�:�g@�F��Z2B"� ӫg&�w��;h�	�ͰXj�)H�1N&]Y>R姥�<��B)��6V�T.�d�+%��
8��Np&��!�P�)�Fާ�� 7&R�OK,��ݗ&r�!.i#h�_ q�A�D�WĀ%�S��?����zx��<�m8�حpH��АNո����{�q�(�$L�A��P*��N��1$l���̀"��cd�,d�8r�;�H�Y*Xqe��PA7P�59�r�Rqo�'�Ü�R ֐
m��b4�Z�/g�d4����f��l���3��2F��l�
0a� l�Ԅz�gը-̐��s�s�Fj�1�4MRƔ�uJ�h�I(ۧ9D�v�X��Um*a+�Y�Ds�*I��֨XB؄�D�zli� ��,�pO
�ȹ�Q���R��5U��Wc�tb<(I�����R�U�5.����rK�'r�Wk��] ��m�Z��W�VȶrB	ig��������H�
EH �