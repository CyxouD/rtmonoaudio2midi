BZh91AY&SYcD�( �_�Px����߰����P�97:�A$�&�Bm4�)��M���'����1���?@
* @� d2h  OP�T�@h4d     s F	�0M`�L$HM�LI�4�OS#�h��SF�i�$��i$�bD�BD$ � }g�~�K���\�ʰl�MC�'.��a�.ch��E�/k_�Ӟ� ��+ڕP#�t��ꛅe�Z���k̀��`���� �!���d/�ae���B��Ɏ;,0�C,̌�̵��*lA�Q��!%u0��+���힣��z`$�0���nx���i��~m6�r\��p@��rQ$Д\��ioH,�jfoFDS҈��w�-,�%j��!�v�Zg�:`LQf�H�P:�5�i���BQ[� �)�rEmn��C�c��e��ECnl�F\4X��m�He{}=i���P1���)��9y�C&BD�0`��ǌ�EdRʏ�B���96U5zTus)�3�F��������#ThG��!��(���:!F]��
Ye��0�+�.Ne��c��~�<�|�	@\ !�ft�)�u��C7'5��d_w��X]챒��S���8���(t2B`Ԇ�hb*L\�.X��pW(VaQ��S�h|-i��3��=w��_[[f���=���|��	������z��N>?���J�i����Z�)�����������I��[L	yH�W'׺#ƍeoYU��?�m�c	jZgg �Cy�����a�!����39tv��9��w:�J�'����GD��/ߎk�cf��~�����v�N�7="8�룾ו$=�\׏9�ݢS�w5�P��߼e�\�cuʍB����s��p0�$�x�DA�&���:_"ӂz��,�f�J(�x	3�%�ɋ�(�.Zx �a�+񋞙�*%U*J��*H�,��s�7�Xe�02����[&�傖���C�i�k��.�z�ʍD ��"q�Z�Ótد��� �k��0�h{dzqu�s���S��vV+��$	vt/�ϒ�3�r�L,=@芐�h$*梡<�Lh��Țu%�BԽ��$"`2��I�3��D�z�u���IAD�D���t�@�.z�{��M�\ %���FZK��^q��o�l�M��ԭ�M.sc�8d3:�$k����*� �ɿm[ЎT����o��'(���;��,���R�*�9�^�I÷i��AۢkOv�h�9`��x�Q<�*J��3�P��;i	�$n�֐	M�J5�C�T���r}�F�%u�ΐх56�Ә�'d%`�4V��NY� j��𩜃+v��P��ay�k����fG��F�'�ӌ�9"8Zi�c��Hf���"�(H1�a� 