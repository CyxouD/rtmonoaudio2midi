BZh91AY&SYukH �_�Px����߰����P�9l ���e�ԕ�Ija2��#%16�#ji��i�FEA�<�&��4M10F&�� `�ȁ	S�P4�����=@�@ ��0`��`ѐ��&��E	�SS1M�F� � h ѠB
;/I�$A$��I!n�� �ﾊL��`�� �P]��?E�Q����D�V�7տn 1��5G����un�6���3�{��RMS��S.��r�����섧��J(�8�	���"2���+��өȣ�RRxDIA{h&��?��0 ̘�W���y���.��i5�/B�]�g�{ג�SY����Y��Ҷ1=˻��DQCq��a�$�U=��<�}':����2�����uNqZ����7,X���x�̓B*�aL	ܸ�`7P*�j�vͮ�u�fq|�yr�J���(Lv��V�kg2���z{NCG���؝��N7[�9�cÂ�m���|>c�I		/�$�@����X���|�^ͣi�n�w�k��Q�����L4�)H�W�D�#�w G����;���H0 ʋ|'4z�"�����+P�n�q�cE����ב�@Y�߃r��+��~,���m�\4kR ;r����F]� ��+�nو�l�tDxѤ��
>$O�.Z�����onX9exn��A� �"�646 ~`��to��r��p؉���L����m�;�F{8.ؼF4�@xK� ��/��l�25�"7	�oMo�!��D�^t�O#5��bgA�}3�VV'Ѫ��	_ݮh�(����UL���$+[Ro^�"�ȕ�Ds��I����7тft�����eY:���-)m��K�� ��Hk�1�Ȅ)�_`�b���1a%�F�R��3��Ai'���@�4f�Pf!����b��5�}J���SH F��35�l������1�\�����Zq4�8���#���t<\`���h05�I��y��(/#�T*��"j>��� 2���8f��3�0�$��Ôu�G�\�c�P'�m�3 �\�H7j�^)c,��^�)R�6{��U��u����I�3�GA�߭*�� =6�!S"�.Z�@��ˊ\y!���%u����4,�R�(X�Ið�I���9�=�M0�91$�U�낞X�Y
G�5,ʫXN�;B�%v^� V�	ݖZ8h�M�
52�E���͢�^��D*J��D�u�y���hZ43�c]�թԜ���p{$�.m�u:�_�6��m�4��5]�L�Z�ܑN$@Z� 