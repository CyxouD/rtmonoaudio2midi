BZh91AY&SY��� �߀px����߰����P�;�`8��f��$�@6@)=�a&�=&��zA�jy5�       �a$ѡ����= ��i�@ �0L@0	�h�h`baD�CS!�d�i2 �����y�
]JA�BΣ�����ᑼ1� '�Q�@�h^�� g &HH��*)�X��;�]��"��p�{�;���-� ����V-(B�33�9~�" xI҄���;3�8�?Cq�lp��䂿EcZA����-�<;�t�i�
�^�`|ك^OA�ŕ������.��՜<��)�­2Ș���ޫj�ɑ~~���N*���ɵlPf6ا�@E�co)�8�"�C*�_�O�Ip7Ռ�`�3X�vd�y���Z�Ӱ�eNn��2ƪ#!�V��i�����lT�6�MzR��S\f�ѴY�d�D�r�x���L��˜m64C�f��'B3��*CY����A�Y��",%UM��nC�@�Z��ľ��bœ�>�79"r���1�Nb�hb͟_�T�	�T�I � �`��t�8rreށ�z٢����ѥ0�@j+5Qj�+�#xt�<KD�0!�Ո���<2��s@ā�8x�0��0�,qkc���O�):���E�Oj럇�Sg��_����Z�>^����j��/,�*ڨ$/��=�"��I	��a���~3%�����ik�������s1�$.��{g�9��!�)���AG�R%<|�4�o��A*zԟ\��9������z��gDҞBʞ优}�@�����H�bzn}�V��ܙ鶙��΂�Y���6gph�jjZ��E�K'%�â�D*A1"/fk��3��8�.���+>W"�>�Y��¢}FOr���ع��UԤ����!TG�p�'8o�:��&I	�N��%
#��)jٯ�)Ց.����›�ո��B����b�3��Մ��W��!F�Xfl^�ϯ@7�#�W��5�����
�L��!z�]K�\����~w%�.	�&	�Q���ۄa��2��6�c�XK���A[~�A���4���΅�#�D��w�`�g;LQ�HY�����z�0���w}�`wP���)�,f��mx��3%��7JNs���\m(�Y�Q8�ZP�������<�#��'����o�k�TP�� ��n�a��֞ͦp�4�Q���i�AN��*��R�Mp�������$*0��k��ʥz/a��\4	+ﲕ�c&��J	���A"V��)}ի�����
��7ݰ��j�FX68=wTt'��8c���Hk�STb��+��/�.�p�!���