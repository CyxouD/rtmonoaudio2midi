BZh91AY&SY��� �߀Px����߰����`�,� 9�UUAT$�L�O#I��S�S�4m(�d�C��T�4)*0       sFLL LFi�#ɀF=Dҧ��#CM h  44d���`F�b0L�`�"h��Oҟ�Pz!����P44d��kq���SR�: ���Y���"���8d����Oh����$N�*)�G��~Gw��^�/j(ǬBRM�vm��i@�����Y�`DC;��ED�t�%�Q�*a�I,�x& h��?t�}ZE�#QBUmf|c��E�mw�Ѯ��ż�m
�� ���Y@
�Πʏw���d!����έZ�]�����mi��PslYl6M��F/����E�C��%3�h"���߁�Zh�A\��
�p����n�#�J��V��g! Z!�zK\�Y`阹r�����Յ;�Y8��K��5cP��f�^���"��'�syн'�jLj2fvӾ��&j����Nͨ��Us��V
�C��@�@^M�Z�/S�����U�Tn#
7�������.
iN���Vi�*a��!A�U�>�-c,Ž�T�o�͍$����azTcR�PC:�t�U��&����n�ڱ�Q3R�[��[��U�H-&�W9�dڧ���Z1*X�f�d��͜=x��Z  @r  ���'N��W0�f�sz["�����d�cV9�AC�����,��������4D���t���l�G/��pBE@��bƿ�wt�̜���Nn��ܸ�����������f��:~�_�ҹ~�^�E�SԦ�#�ћ���ʺ/�UP�i�G΂<1�~14k+z�#��H���5	γu[���Hx�M�$���)	)��n;g�ar"�>)�����8Ic�+�׹zj��4��?�}P縗7ư�K)�!�<�w_V@�זvs�>"S�v�%'��d�-�t���d�6<��}�q-@4"�TW`��o*��b���V�aQ��#�Є9�i�C��?1����Bק�Vd�jc]��ϝ6��c��<s���	{Ӄx��P�1�B�F���0!�`����.9���3�
S��c���dگ�Nh�i�F��fk��G� ���}�F��1�<8�Xj`@�B�Ҹ.@gr55��s=ȀV6@�D�2D�[�F3�\K��A�����C#F̠�}'fJl��ɶv�EX(��<s7��(���y�y;wI�DN�Dn�IY��C�
�z��ΰ����+f��mW����gd�#��q�)=�BڣW�@���Y�ߐ^�C�xP�t��mG-ƥrU�d����6�@�<z�p�3�6
����
S�2��t��%������kt�M�1���r��N�ٔo%�<8m�`ur���:s���E��>jŻ"x^�jjC�����7JN\N|�?�&�D�99g=>-Of6o{�5�d�X;��W�.�p�!�?��