BZh91AY&SYmS�w �߀px����߰����`}|�x �8�YQ�:a$�4��4G���FS#��A���j��@J��!� hd�4d  � �`�2��H�&���=@h��     JI�=OP��h=��  2Bi4$�zj1�2zi?T��@4M7��~@5���6�2�?�)��N�m!d A��9z������'(�����w����I$��u)$���&����5����	f�/� ��cr�JmL��']lq��UT!!��[�m�nl�����Ln�(*Q�J[sa�X��` �M,�?T�6��eɍ��lN�����sϯ�C\�iM�t[��앒���K)�B���x��M�
�O��d��K�)���]�-��b��i���*��1� Z��z�V�c֞��7��7QN\5T�ZSu�b�,*4�� ��)�]m�K9�j`n�1fD@#M���lx�̊D��~� �&�DC�b�4�],���0�d��bTL�݉��2�>��l��c�3�i���+'D��\i.N�ԭ��hÀ�v⩜S�Tdt�lM?K�؃Z
z�q��� �6ËX��誇cKIt��UL5܇�"�����g*1����`�R ��$u�"���)uF�;�kj�@���ot�܈]9|Z��^���5Nҙ�E����̞5��Q�V1Z����ԂXaU�Tr²�z� mUu���+l��*�/ (.I.Dn��w99�D?ϓ��}������m��0  �W�p)h�K���3�V�^d��"��}��&*�$CB0���x�~���DxZ���y@��^g�;�d��q�y�LA	%F������������n��=�����Ѫ���/�����{�?/�������O;���JI$�������u� ���Y�a���q4hQ�)���1  ;�?��hv�G����:��$��������ל[���TA)~J����,=l��������j��%��� �{5�Rws!0�H
X�Cv�M!�[$�}�r�%('v_m�}�|�v۠�����$Ӯ���ވ�-�R%Q_��[^����&6O)���0E�l�I�B͵LV���W$b�{"�m�'r���|�Wq�ǫ�>X��:z��XP@ /v��zܡr3�f;�z6���?�����]��ȡ�B_2&Cm������57	$�i��a�����tz�9�r���c�\�$)%{{@sRtO&O<ꖤ�lOL&J�ww��~�D͊�]�-��C�;,�ӻ���6l�}��,)�un��a�Y��[F����� �u�>�A���'BlI$�RI,�Z��=EE�N��ח�Tr;<b�h+/�<������2�G	�]��2cI �Mb�~��q �4�.{T��Rnٔf�%@�% �1�;�UD�s`x���7dI������[,�+��ez�V7o�$<����4U]b����+�g`sB��Q�h*֒�4�m��HxZ����/4a}����i	��e����NF���t  ��w+���G��dm_�E��P�E*�ܑN$T���