BZh91AY&SYbl�� m_�Px����߰����`
?97n   �RR�BI��MLi252yh�i�i�&� �?
U       ѓ �`A��2`�S�?$M0b``��&�4d���`F�b0L�`�42e#���CI��<S������z�jc��<����D �B�� ���(��_�"@��r�Y�`�	 C��R ^t 1"�6��.a{]��?�V:D�T��bY�A{�A���&�mn8�f��E����%�f˖L̑��lm
R��Z��B��.�K
I����n	LJ1�ȉ*���Ofjt���òvDf4i��dЂB�]CD�H艵9m�d����yU���!:_�X]���O"ҡ
��@C��ũ�DN�Z.�|d�w����H&.��9��N& ��M�����.�~�H�0�J�ͥ���i�T����3���X\20f�&&� F}x�
��bEG��,#/ۂ0@r�DB�nmȩ��$簜TǑ#����u���X�oMű-P����r4�XJ��G4{���^|@�%���,�&Ql�f�j�8�E�Є��L\ޯ �QhI����y�3J��~�d���E0��e�Di\`���$��Ze������O�es@�$�q�|ğ�e��=�w�����vha�T�$�
h�e�Ә7|4��L�w w/0�5������慘/���yQ�R�%s��d�f�A�U>#:߃��Ҝi&�$����̥��<�˅�|v���`�2����/�pEƨ��_&,FE�i�ds�*�Qz������%7�4��Ou�UF��N�̧P:����(a��P��~`J�\�'��TUY	���}�ӳq�b&3&����ّ�N���/�Wm̧�.w���᭨������<w�*F�d'[3w;���#�z%E��ɘ�d\�A��v��3ۮ|ڜz!T�Ag�'6+�xH˶������f�{���j*&D���P�(��.�<.n&WtR�7��"��f�k�dft8y��r����4��&��^�[9P,v�����w���B�115w3���o�u�?v�۾�]sV~�j����p�eU����6�f���1lv,�T	]L���;�uoX���wN�u���|`4��j݈{�:c��Ta�����t��\/T��<�
�FpWEƨ^U��k��BdY0���3V׭G&��A-�q����U�kl�=DR7�*N��J�wc:���������N<���-E(���ƿ�{xaX�/�T�d�6X�����P  �� ��t)��)r��Ub���fK;lL��^���a(E� 	c�� v��b*����%�"� ���ƈ;���Ʌ�گ���� d̘��v��Q�%ϗ>j>K�6�W����~>������\W���6ĳ��*B@u���/"wdI Nc�H�o��c��ac֪����1�� 2����,�`�B�E���ؐ�B��D��{j�z)J������qA����5���:��	 ���:4����	���|��e��$�,�]yY��JT'p���+%��e�"�ը���;<�@��[��X��ZR:�2���u��f��J��$ 3�!�鋪#�\�Z0�'͙�Lד!esQT�Na �{�^�;���q��S$��86G��c�ɜ��@��VH.����P��Ri���T�_�)�� +��61뗙��ƤN{+��,�$�3SB@���^ sB6����70�#�TX���YD_�+�4ƌ$�b��NM @@���ډ@R�)�3��F�QY�T�h��&�͎ˉp� !T�j�&ǆҔ`$ h 5l"�n��L�MC��|��8^o��ɽqv�9��j��6��Ga���ic �z����[��P6� ʝ�|��l�ɛ~����ŭ�XXe �3ۙJ�E���ʚ�l�a����+_�"��|�V�4� L��U��"@L$ B��&�R�0���-�
뫕A�=SlGJC��@uH�.�$��4�z(���عb�M�HZ���_�ӥ��BH �fGq��,K�׳=�	�i�#�����H�
M��