BZh91AY&SYYAj J_�Px����߰����`O�[p��U@��QP�Di��4O�S�OML�Q�4���=F���R �     1$$4 �C�    j��@  2h�  ���&L�20�&�db``$&�O'��CAG����� =G�z�АO�$�$H�����$�S�?����b�*��E� jz�l��Ą^0E�m�!�U��u��-/��{��G�	3���5��V��II�E-9r��b�I2h�H.�T�@S`��n��_$�&\1 ��n�}��"C/f#��\���durH@Ye��\'0���E0��?��=��ͮ����\��� i�/_4:�����6Z&l��D�\Nf�����dA��V��o" 4B��(֑���L�	'���y���p+����UZ�K3S�;�U��c)h,����[%�#pn��
��A�ܢ�d* ���QhCB+0a0�7x��d���$�F�%(���`�#���m��5����m�8b��lJ"��J��=.C�+dg5@��aKL+�VⲦF��fJ��,�l�O�I�i��wл�ؐw��#[�c�0C�62��-�����Ð�2�~�3�(A �$�@( �X*.:��H����\��J�Ҳ�Ю&�DC1��
W�х�V*0������C1���0{���*�Z�<�Y����j�����3w��y�UN���c���産�ˣ�_��fa�Iu1軑Z�|�{zziD}䲺d>�%٣��Q�KAC�y���m����
U9�n
��~D.�Z�������u?ڜ�u� �������s$0�J�W��������Ƿ1�Ѩ�9d��k� ����͍�([._u�#��J٨ߍk)\۰ˮ�:˂S�P�gd�g�88ؤ�4�F��A�Nt�F�}X��yy��TiHXl�3;�����FCe���ēz�_r�Mz� ���\܈������d@�sP��8��F�T�U� �:�;bK�� �2f/dEN�S0�O���%�һ5�g
a���=d��n}�"Wxo�����tb��^li!� ��]�i�=���s�"ax��P�pjM�P������N�W4!&��\���j�J�DB,��ZT�[�����&F�o  @�2�?GtA5w_1��V��d�d0�MQ�P���|M<�_�J��67C���p�u+�G	�7�[����@���kL=�-z�5� r�&�c�26`��U�Y�4��V�F2`A�pn)0��y�f�l������m�sU�������Y���Щya��ʀ��2�8��r���A��X��nu^���	�rZ�!� �)���\He���opv{K2UV�8�6��MF��J�dx�kً���2G]�ݸ����)��:P