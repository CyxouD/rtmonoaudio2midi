BZh91AY&SY��^� �_�Px����߰����P�[u�q]���HI �4ѦShCCI��Ce�mC�yA�~���$ �      H�"S�&OS ��i�@��@4�� � �`�2��H�4d��$�#M  D~��@U�@2	?��_�$�~6Te�6ڄ�P���e"�$ ��ch�a"�2k�uv���RZ%;o���t��:�v��f�eIi ��E
IJJ<�v ٓl��s5BFu��1��
ւF>CQz��L�̃4C�@ �!
�wPf��zn�d$��fM��N8��������C������Х���;�kN>�i�W�1y�dqBAx�N��%#���ōfSE���ژ�A��چ�jaW���1�$R�f8��<�&у�6;A�H�DM�0A��D	�'eM��KRm; q�S;Q֛�mR���B�I,E�h{vУ3+�ɶ�9KZ.b5�F��3�a����R�wUW�-1���l�g��ڭ*Qp�Y�V�)�E�&�DI������²��+r-QB�$h�a���X��9Zgg�n�I��66�m��$�M���:�Kջ�UzVy",�g,Ejk]7�l"\�H�F�:(	b���"�I4��.�����`�y��v�BM�UN+k~��J~�S�O]�[��?%�/���B\�P*������?��c1�¿ڝ:�,��{UIy[���?�V}"I1L���@��b={����5=m���;>�,f0J�+4�������8�BKd6p����r�l�WfDR��L��ˉ�:?�К�����b�D���҄�^��l��:5GfR0�)\~]&�h&�}�j�%�i����e���}�󞔫Pג�L�In0�KFC "�A�L-&t���TGc��00������虥�yMW���}D���+{*�/�}	+x,D�G�tulҘI'�b��{AkO�Mz��uj!�$��THZy
M$ �w9,mA�dֳ�}��k��W0�0ֽ�?� ݑ�;y�L���9�X�pTk`H2BK��q�"���m�a��T\��������;�Lh���D�M��&��	@������T�E�����ĔrL�e��뜰$��A۸�	���ք�ޒtXh3
�V�����U�#w��'����9���C0s��#I�'q,e�	'���G
d��k�	'.y�'����K*1�liV�Pp��pf�N���: �Y���,�0U��?H)�EAP�M5ju��&)&2�ƙ	)2Q���g_B̌̅8�j
�4�+�ݮ��"C�7�$V��ڗ��m� ]Wʖr�Ě�:��~s\H	%X̏�ؗ���r��2d����4x����)�n���