BZh91AY&SY�)Z )߀Px����߰����P��.�#�aY5�H��	�I10���)��='�zOPi�51�I�F�i�   � $$!MdMA��  4��101��&"QM�x��I��4P�hPy�(6�����z�����:�$�T�0l��5������-	��K@�>=�{go ��Ym%3��v{e�xS��+C���q0�c��J\�x�Pr��������[�uZ�C6����B�=��Cfv5=�~D�O*I!c5�L׈p[��vx�`)#n��x���98A�|ͼ����<�t{,�:��q����BK���$�1�n](ɜ�1�jv��KeE��v�Dj(�)����ٔ��h+fM���kzw,�A�vT��L�V�ᜈ�̤2J e@
��9�p6�\T�Fo*�`"E���O
���=Z�;���!͚���HJ#X��M��:��K�ZL�&	]��]�a*��
&Xn2��Yv%8�;K�I����k%ʉؓ�:}����������l!
Ǔ������+��r�$�)�r^�y4d=lхdM��Sc)g���F̘��#	+\�%s�X$0M��k��$Yc��/�r��u�Ս�G���hKo�Ag�������~>�ȼ�ʼ�:�[�V�0H�o���Ю��S����O�%|>ߍ���-���A���˙��Hα�w �&�p��,�}��H�F�n/�(������kw����B�!��a�J>�ƛ��s/Q�{����"^"�Y���p��yw&��N�Av�|R �T�祝�W	N)�m��
���QVS��F���,x�lL�� $5SJ��k�Fšm�`ئ��9qu�)+�-�&`mr;�A�k������ejJ��|"��8�[D�p�T�02!��A`�4p�R�V���zH�Zl&��F&��{��6�����Յ��H���36l�] �hr袹�c++�*4�p��P2�w��oJ�3$�	rHvA�E9ҩ#�32'�"�D+d	8��^[e�����3�ݺF��Yd��eVP��)L�y/9�	\&������qB1�`���IV�K��g
������3����X̓�lû!�:VH�A3����«4 )5g�	�²�ì;�5�n�l{D��Y��jW��cZ����b��|��#@;�
������y��mխq����X�5Dk��@��cw����9],Ӄ�e
5�(h$JU��:�UV�ǜ��p�E"��^	{+��9<q^��˷6�W����7np�.��6*$����1��$p�~���]��BB�h