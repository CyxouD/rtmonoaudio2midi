BZh91AY&SY"�� �_�Px����߰����P�8� ��43j$�L����)�I��4zj�56Bi�H @     $$MO(OP= �� �101��&"Q����mG�zhڧ�=M  ��6(���En�� )D� 8TZo=��Q������H	h�@�� �` b@K�"t@�R�GnO'Nlz��ڻ6`�~>�A�w��w�{�w�o�JCm�5m�GѿU��c�e쥵K������kcu�*�X���^�s�Ŧ���YE3Mj���%�5PV�m� �>~ �w��o�
20w���V��Xr��z^��N=�:����xl��3��l� ��QA�7SM���C�N��"F�����M��A���½F'��l^`ql��B0�t-���A])�)�i��6���3,i)�Yu�\�pX��՚���yX���n��ʶv�Y�Z;���E4�-P�GGv�\ �Yhc��|�b�S���/��{��Z��Y�����5����#�5yG܃Rzo�{��d��������ܜ�M�66�����!Yx�Ur�/�-z�&L�m��9��f�ITF2l`1��mbW�1����y�	�͂E�r���X&�(�_�c��2E��sc�~t��I�g=9p�{�l�o�HO_�r߇���:?�O-�L����$��p�b����m��~%�b�e��\J��%�w��#�#�qt�|�ӻ��ñ�sbH������	�"^"H(�(��~��k���o�Z2"IW�'��#�<jëW���@x�$)���ƻ��{'� �-"�n�n�"Dg��s3����"�����]L��y(O3�L�7�~�n���F!uX�Q��T�R��sL�@�ny܎�V�JL�$&��Z�LcY>�"� �a�����L�
��T��]nsjJ~*R�[�C*5�����[kEUhUh��ٜ�:�i@]�u��3��H�1{h�"B�zq�@$)[��a���}��z�<+��+)�cm�+f�B`���.``���l96փ�!`������0Ċ)%"��ъ&���V� &�Սe�����3tG�4j�]V*����Γ��\*4m
r�^ӗ�:⎑GV��9j�`(퍻�~��-��o�A�ػ��}{F`M�dt�[�(��<��0���Ü2j��N<~��/��ѺV,R�:��b 8�sm# 	��!��j�YY���S�*t�!VZC}w�)E�;�
�J����$*�HUa����0��h�,0���]u����p�E"��و�r�������c:��*�MQѧ!�[��)!\3#�ҥ6)�T��t�L�5q�����H�
B� 