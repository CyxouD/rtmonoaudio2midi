BZh91AY&SYoF� �߀Px����߰����P��[�8b�-K�0I" 	���ȣ�CѨ�SM������a%@��P @  "	4ҞI�i�C�= �4hh 2hhɉ�	���0 �`�0��FI艴��M�  &
���*��)!�@;f,�'��Đ��+)e�6�HMC�YH�t� �"�P��C��vo�L�[6p���p�Mo	�˳S\eٚ�r�"_�z��9�FP���e�u�X��y�%(�[.�3��蘊�]�D]�-�'��$��{������r�����5�w����(<E8�:1+���DR�xXX�[��!�����#"b�EF��� �#c#2�!��" H�ep4E�KL�"#!����]t�F&�p�,`�,�^u]SEj���f
]�bDU����[3�&�KlۭM6F�g�����
��(a�S�
!p��"PfeK�XwS!�V�l"�$E�Y�"��ÎZ[҅K�9�fbu�c�SEeH���p<��'��|��PA6��T�IK������툳%������'4E!��8ir4�>p4�(<Y�"�!1nac(7R腙���(j�	$6��<=]������,��#:?u�;�����z�/���I<�eS�y�2�e�H�eZ����'�bi��,_��y5���/����(���d+f.,�4tnѷ�=G/�$m���B�~�By_޽�E�J,�y�I:�U�l����_��K�c�zqT�)!Iؖ�-�P՚!��ޚ�����2��+��(����s�{��Ya�h�}.�ٚU�C�����HD0�
�@�Jd▔�N��L� �:�2�9YW5FS�Y�,�[�b�C,�g���&"�U�x�I
R��.E�x9��� Y͐m�L4��5ٓfZ��7qx�	�b@[,�Jh�4
�rH�-�5� �q��G�I
��0��y���9��c�mc	�N	L�$"���􁌓�6��X���������Qz*�i��4N���j}��H� ʘ)N���f
��*��B\�!�D�y�r� JB;ۮ	���jE�!hI
���
 �T!��O����;*z
��݀����3�G~��{�f]>:l�`�Hv��=�7[U�_��V��<���\���@W"Z��ʫ	T?Htۘ�H��Ñ���(h+���7��HXkτej�|*6gª���Zc��H���q�u����$���Z�aR�g#O �w�,D��Sq*5#����P ���4(cbN6Z�c9"�L�}�r��w$S�	�4i�