BZh91AY&SYI`x �_�Px����߰����P��nƵ�#-\ل��d��ji�42z�4d=M2d��5(�yF�F� �Ѐ  H��S�C dOP�=M�4 ڟ�=C�2b`b0#L1&L0H�b4�Q&���OS&�i� 4 	I\�(s)J��7H�t�%��,��0l��j~t* ]4 �"lm�A�M��m�Z�3�!�)�~�����a�r�+�T���2a�h�UD����cnM9�#��2�y�Ǝ8�#+�@������=�1	��P�Rv�*.�Cd��g��L ��O<����5sB��i�*�q���F�����C�p�։ǽ�q^�:5��ހ"R�)K?��B��J�=�`akk�»��_[WE���#���aA�2�%Ю!��+\��I���B�Zڐ����̌a�k�ݠU��Y����<��/J�	b��L �I{=����K�ĸΖW���<q�α!�vi�������6�l@A���S�J^�|VWէ�"�K5DZ�k�R���l��3T_L���B�"� ��a%�M�)�(0��u�( �M.*k{�(��G|ث��\���c㣷!O燫�w�ò�dXU�M�9ba�J���Y�χ�1$�}t@��96��t�<���U�}]Fә��,f5$U������@n!z�r46 6�`7Na<�+�_̲X����9��9W�=�G��g&{�8�ڐ��@���\��ǐ�Y�Sʘk�"|B���h�Hg��%���v�"R�vڣ��T��yl%c|��wr��9��2/#���8� ӵ��[�]�`�Tl06�$J" q'�ɖ��Ae؃!��wo�)��I�ƪ�K�@T����@�?���;.L�zprX�$��Ov�����9䞖jI݋QA��A1�ce-w̳�N�X���1��D^���t�G��~�j�5f��^�κ@���j�S�pT|��h3�)%"��Lh�HdRw��I"�쿪H��0R�6B;�H�X*W����!ܢY��^�� !H!�%�x'�fD�� 4�=�x�oڮ�d�����!�#�{������l����j��#�l;uي����ǔ�2.�� �D�ܳ�s��`2�
�����v��bd�;^���\:'6L�[RP4�9=oKN�R�Df��e�B�5�ĩ@%
e�����dh@�wV�7�4�W�B�ȅ�k.H����/UPl� c��灜�^����IP�]i�K��	����h�/z�r9�2F��n�1�rE8P�I`x