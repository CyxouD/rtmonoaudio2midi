BZh91AY&SYEh�� q_�Px���������P�W-���"��B2	��<�0�M1OSz��L�Q��5� � LF�0bhi�L0�ȦF�@h@A�   �A�ɓ&F�L�LD�z�z�4<��mOH� @��(�,riHJ�H��"@d�J��t�?��e,�� ��0�\M��Dh���v0�H�
5�z��-����nQ��@K�撻�+(�z-pl�+�Ik����$��uNj$�
9f߄�*�$��܄�Iƚ2Da��I�D����ja!+����8m�����!6:;��ѣ�������wG�ɕ{�O��~�C~�ls�)���ֱ9�Ag&S�=g2��5�*�w�j���a#CI�g*s�RTU�|��g�
ѤΉ�:BL�5�`E0�Q+B�/z���`�V�٨��5R6������`�R�
*�v�F���$ҍK�J�%�P
�r`�A�G�vlP���-k��*��1����|"*Cb�|EN-���	��J�%&�ىޭ1aE��X*ӫ0���~���i$$$��$��M��Q;Ɉ�o�e���ݑ(���Ye��`Hͬ�ϣ0���E ��]�<*�fqS�� �U�ś���\�x�!�I�����3a�z�d�>ysJ��d]����/���׏�f%�ř�ub_�͊����w������l�,�_ʲ���n���������W�|�(�elԄ.Eɳ/xw���̂�*�����n��N���Y�D���W��z���	W��N���Z��g���K��]x�+P�9���c��T��[��8�������T���8��}4:r����Qju��x�2H44�(k�Z�C��`u�6<�R�U4�N7��3	��,݂0'w��E7��lfVR���1_(j�(�P�����q2�
RPW*���^�^�A!�h%�E�\P^�Nb�9),��G0̏��H��,�cV���;��~9��B6q�U��f�r�!a�i k/G�q����x6�N���������H���M��ƋЌ�b��  MS�|�H���p�pU#0�R���EH@�jfw5ĬB�a����^b������*h:ys�
[%vڃ������Cw�3�Ԑ\�0���ٴl8,�#��=gAݷ+$�O��t#�2.����PUt���q>[�2�5Ujʕ�%YA��%\ٯ*�B@�C۬�,Zr� 0ӜG2�'+P�$��h���H.e��X!Q�W�	7�ł0df@�9�0��:,��!J	���H����/5zۼ��X�\l��Y<�F�Mz�	! �<M*���Y�E��QH��H�|:��w$S�	V��