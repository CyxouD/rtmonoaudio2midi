BZh91AY&SYh��� 
�߀Px����߰����`	��(  #��L� $�F��$�$�����OQ�Pf��mB)�@T� 2 0&�@ sbh0�2d��`�i���!�HD�HѠ�4h �  h����&L�20�&�db``) E?J4f��=C�d�4 ���R����"�+QQ(����Y��|_� �����_@K�� S��Ո+�-���"���>/nj�	l���H1��Z9b��h�?< �s� ��ä)uUU%$�d*Khd%������RB��p��G8���w�P"1:,��Vu]n@b���W�A^M��\��J�ٍB�πq۳��ཀ����J�˰���x����i�ːw;�e���q�}��Ǟ�N���SZ�wp���Y��2*��Xb��A(&�N�́�I�U�0�)#��\�b�l���^�d<:Y)���[�U�Q�y�]Q"��%�އκU|Bst�:�Ҕ$R����q5���Sq!��3r��ܘ��1&{�1a��C]�9 �6b�4��k�3�u�CFa��k�� �W�쉲���O�,��~DS�##�|��4x�NG���<:�TC�ZH(�k.@n�Z��[h�ѓ�맄u0G�GУ��xCÅ e�oD���=��*_�3늑��M$Drk������@T��	Rh��싮��d���JS�uj�p<e������@�RĘ�=U��0w�!�DunR��v\�1&�ˠ3�y!�֤�I+&]��uO]U�mT� UWa�r,T�I�CJ]�d��2�����Ա#��P뱲�u`�:{eE�Œ�`qO��&*�6%���wss9�%�'9�V���05��]�>P�Z%�ET���ś޽��c5㪮�(7)�0�6:Ds6g�bF�d_e���P��פP��$bq�</��lX��R�^���S����X*�[�����勾�ڷ�ќ��LEFf�3\ω��4�in��s�H9	,5G)ߪi9-��U�qT �/F�w+6z&k���S�n@�v�� ��9���SQ[�H�}Ǹ��{uqn��j:��G)FH{ws5$�i)Y��e��t�?�J6��o���g�̱�?^�^/9�m���Km���P�e��*�)/Gw��I�)�2c	fЖ.V�#Mdhĕ�	1���-��1ZA=)h �|�.3��+�v(�sl��4�L�+Ƶ���3���5�ק=�'�uSsx}!�3��%�~���j������ F��Z�����������3gB����D�ʂ][��� 4�,��_��9�u��d�	hZ6_����ï�FC0 K�:g[�D֝-��h�J}�D��Wu�Q�M���/�Ɲh��@�*x%��V��OB5�"�1V���X�^ꗍl���%8�涚a
�����3L��4$���:w�;"�$ b�Q�[BATN (w�hڸ_f��`ug,,��*�[���Xl2{{DȐ�7-���A�n86��|���Y�8�M]��N��zj�A��*(N%�F*�xq���ėƠ�X�L�[J�q����b��ۢB՚�XJ�%+40�0�A��7�C®�c�ffTȠ�  ���0Q7��M�L��XbN0�%�H�EIvk
��L���̭Z%�{s�(E��*N;��H�Z+O90���,!Y)L�y�1h�-�
��^���vS�.� �:Ҕ;4�;#f���;�g'��+i�L�>I[�Sx�s��~%��@Ag{DK�g/ f�$�[���N��2���ŝ+C���b 8�E���@�y��%Vٰ[�w"���
����T��V��d
�\�i	T��*-���i�I���\4J��:�5Vڇ�� :7H�ѵ`X��N�r�4G �F˲(�R��Ә�'(�V�#�4�R����c���Y2G�ՀW���"�(H4q���