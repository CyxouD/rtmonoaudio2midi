BZh91AY&SY��� �_�Px����������P�މ��2�6�$� SOSM����7��M���@j�4�
P� C@  BD��e4�22mM  � h�S  4  4�@  EhF�)�5OL@�i4� ��4�� �@���0J$��P1���_��s䩘`�# $�a��- �6��)ch��"�k�:�ך̠%�)��S?���|޾�ђ�&�\,N�y��Qӵ�:�ub�e�b�����h�ki�P��X��6���C�<�C4�!�+�i�k�T�[�BJ�+��+�`pӿ�w�M0ll�,����9vw�[��P]��[8�&��hR�! K���imٲ�g�Ĵ\��Y�`��*2���r̶��lX���jf�L��Ԗ�M���\,�y4�CR�b���i�[�u�BX8lβ&���d�j0���T�a�)e�ibC���@/�a ��W2)�(��3�nm]g�Q�4E����n�m�H8�M��Fh��lJ2�	�*�13m�дuM�8;rZ��Ӊ��qve�([;��k�:�Aa�֥ϧ����f������`�%V[[�Ȥ�NK��2��e3f
�d��1d:��7!��-z4���T�	1r�����5ś&��^�i���#����N�,��=ܧ�sF��������ϛ7׻�E,)�כ"U�}
`�O�����$	nqM$�Q!%��㌧	B���)��:;f\٭ZV���* � �Q0���	~� fr��&����v��D�O�9��r�7AC������3r�:ɽ�%	nb�������H�(���U
A�{��/�9��%4���^��S\WǍ�����D>lr_q��A��)�FcB	�4�v�tmZ��@�&gwQq�v�L�Hf�1d�z(+bvr9�҂N�R_������Z!�z�ۥ0h�T��jR�7S��BC��K�a��L>}ef%����3+��$G"�V�q�*-���;��O;������-u1��c�s��@h,v��.�<O����8����A��H�JU$�cD�Cvb��Jք�}���� ˙�N=���f-
�]V*���sع��  I�Pv1��H�+�KN�(6��X)0��iC��͉���}��OAS6G9��t���\�����{�J/a�I�Ͼ�@�i���Ϩ-�NR�A�7���U�.ЭJ��5�(c$lϰ�	�f�/�������8H�6�r��B(�Rr�( a=m� %[*r��z�W"�AF�Qȥ]u��/�]���	$�r�X�#D�]V8 »�V��r2�_{��"���2�b��3���HŦ����=�g�]��BB�Ӿt