BZh91AY&SY	�� h߀px����߰����PM�n�\d���	$���d���h���i��Hi�CM��M�I�z�����  �   $$�Ѥ'��d�dh2 i��L�i�����a�0  �ML��iOԌ�	���~�@h F�T�PHzC��28I����!ty�Vfl��>��_� ��Q��ias\���|+�B�>�3��������G��K�mC�H*D�J�?�:1cu�V��P�����68��ё�A�4hR�7� �tp��)��������nK������	���7j_V|?�Dҵ�:+&�>�t�U��{���0�0�S���(H��r\mc,2��"_e���:��=�,�xUi%��
04) ��R3���|R(9+�\Sٖ��$4��q6��8w�%�-�a�n��6FLk�1���i�����˳�������m���(B����).OWn兮�ԗ���K��2����62��C\5nl�SJ�,��Bip��eBv*\� �E#��O@�9#C�Ҿz�!S�{�'�qK�݂��'c��]���޻���B����K��#���S�P�����MV����DS��M�������O�n�ܿ�)f.HXU���i[�7\��hd6!~�`7��'���kZ��d�q��ŵE����<�G-Zq޽-ʀ��B��_�f2P3�Y:NT���dI�z*|�+`�q3���(=;~�p��2ͺi׆ن����w���[A�k��0Q$4�s��V�l�@�*eGl�՘��N)E�4`��B����A��r�9Bo�/�Uj��b!T����-Q�}y����|�V�h��%����?�
$�N@,9I�#ެ�Fe����"�`����Qυ�a��&�8A�L�d��nŞ�w��aS;@�"�z�$�'����đ`T{A��h8��L���0�i,�b�A�{0�P� ˌʓ��lF���2�xIr�R��B�R���Z���:�W,5��#E��~T7�T'���F��a8k����UAA[��l����YG$P�y5�l1�O��P�ɐ�/n��p���Hl�%�D�س�2��mHj�I`62ĤKObɄ������8'n���ݘ�t�ဗZ$��~u���á}��Q3��
WvjB�HQ�Mu�\����T��zD����*�#�/�>S3�g�!%*U"�L���*��Z���~l�&c��$\ɒ3P��o���)��MVp