BZh91AY&SY�k �_�Px����߰����P�9l⣸���ւ�"y��4�5=	�'��M6Ha4h��3DbT  4     �D!Hi�L�h�=&�P  Ѡ���&L�20�&�db``$L@��ب�Щ��=A�2�<I�� �0� ��%B�x��N���G��ꢛ*��E��0�}���HXF6�&�(��wm\|���4�zT�s1�J�6�,�^&)�*��B���q��.�&r��j�1��~O�IB���QD������
����1 Ȟ�Yҕ�A�Q��	
���!m������df����Ű��Xf��F�6�a��m|E��6�&XC�\�6h�ƒ�H�6��!��Y�iC x�^Ћx��282��õaQVTBSG�9�bЕC:U�L]�lL�k]*�ib1@�B[:,��K2�լ� �,��r��`�����r'7u��:/l��+Z�2E�Q��	'f|H(��;݊*�%#�h֜��*�>�~_1��^��I �������y���*�z��(��3��I.us��M��4QI3�:(�Dt���*eW7\�^©��������#P�-f�v�H�y��^���.�~5���(���|p�<{�M�?|�<�Ny�1��#uyt|��l�!Q@�琹��-�vJ<ih(z�>�Y���u��!���U�6Y���!}(�:46����}�y٧���7js��r�Q�K
�q�^�r�8-���o�/;;s�ME�Ip�\s�L`JdV���vu�FD�Za�eLpy�[BK_#�9�2�G����@J%A����AB�g&�2|�;�G���ȸi\Ԑ!����j��SR� �c)���$��`S�׷�@�˶u>Tq�I��j�0b)(
��vF�ܩ��Lo�MQ��� �/c&8�E{a)�b�`L��W+%�� D�Z�0�X����j�s�עY㥎gNY����	q@���ud#s<���"a���!��I��-cLh��̚t%f$(R�k�!�RN��#K�3#(��v���1�2oQ��2�,�ʠ��썈ځ�#O�<ym5
|��;��˄hq9:�jz
�㳛(���H�9M����64|1���$�]9��|"���G���:������,��ˀ�8��'pD��G��p�˭��1�l�L�m��^bJ�T\�m�
�(q�7��{@�e���<w⨍l�+jʭz��}�>ZĂ�@s&�L���ꕟA!l�.���3i�!
�T�F������0�`�u�_�#1��$cd�����bЦ�.�p�!��(