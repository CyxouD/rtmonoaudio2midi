BZh91AY&SYԥ?& �߀Px����������P�8��#9�,U0�A2	��S�M=��i��zF�mFC�G����E@��  � �`�
d!L�4h�M3P � �&L��L �0L�0�(�Dhh��yM��h ��[��H��)D%3 �k��}� � �(�0k�L�
�[Bo��R���lv��ߨQ�c^��g�
u����x�Gn�)���I��i���ܟ��s�F����3c��,���� �FP��ӱ��w(VÒA�]��7x�sL$&``����;m��8��.d�5��uv�.�� ����28yI��iW@��v����Ad�B(av�����ϙ��"��h�2Y�a%�-9c8�t�K~F��"�*-��h��'IV ^j���.�#79&��@�XPLC�5˳�0"�f���QIRb���څ�cr�*fV*�T�f��]� 0��-CęQVs��"0��!�("Rn��/��!�]7�V�,��J(�8�Q�Z����N���������H$x[m�$( �l�S̉K��ׂ�VV���Y�rf�
m�0�r��@�Y0��A�I��LEĄ��0���N��f��	��Qs2f�b�,k����]��U]:8��x/����x�>?�����S����Ai�_�7<��{iҦ$/,����*�䐩��-���#�_���F��౯�;�Λ\�HY�lm��7�{]B�ld3	�s0�]�kvǝf�J{���Y7Gѕ�oԹ�4i@z��	
D��9-&VN�1zDt��v���ܯ��43���%8'sY)=�wM]���ʩj��[l�P=�
XKF#��8��i�ɝA\0X�����0��AnX0a��y��� �G��c�����r��w��By.���`!Q����=`�4k��E����Ҟ���~|J�� �w�1��n��e��F� HQ�3�s�Y�g�������c���ȮpV^�@b$|}Ǽ�L����Y)@���ER�aI�Q;CLh�����N- S뾢DP��Jp��80H�X�N�+Ĩ"�K-f�1��	h��P�>k���t�G@��tA�_h���z�zΰ홯�ٕ�Aas��]͈��6H�9�S�U�)��a^�#�0�p�����y�}����/�Բ�@rfuWXDUd���)P��	�NөLk�q60�C�
S�"��|c;����Bc�Jr5G4
5Ѧ�L��S%��MDP������׎�Ǆ�pj �E�_r^�ūa4.�3�c��$�ST��i���HY��^�&'雎[5��o��85G/+7M��]��BCR���