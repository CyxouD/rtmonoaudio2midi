BZh91AY&SY��
� a_�Px����߰����`_�n G{�E(HH@A6���Ч��H�A�di�jy	�J��      ��2yOD4h��ɣM&�Jz��OS#M4f����L�M4 ��2b`b0#L1&L0H��M2�U?#��?E<M5��h���4�.�D��؀EX�4$%I��{HJ=�}D ���lSeX6��C�_FN=&E�X����EZ�˧���� �=m׬{���7�qţ��I;5U���"�

)���m�������x�ዹ.���~�ꕶV�P����Fu�4IBg�-'i+����cn�S) ��_�l�Gv���9�{���ͽaO�؛D�6�W~I;�pf����N朳�W�ڼ����nL	����	#I��O����$ N	
8�d�Y�n����c%���Z�f/��
��X���E�5Y�i�R�D��}$�`w��gc��Z�X�N�BH�n�s�0�;�X��� ��&��5��� �����%
�]�6�@ʫ!#Q�ie����Bt�Ͷ"�(E�(� ��Ywvq��
�2��|�e:�DPt`�:�20��Y���m�M��+Cv��	���Q����8V��}b�u�v�n��n�|�iQEx�U ��JˏLV�Qx1���)5L��#��A�@FLA#D�2&�����~,E�n�bg"]�(_c���0�akT�2gK Ў <Hv�Ѓ|2���1nn.0�r�0��D�����,��.+�U��
7S�LB������WgH@�UP�i�/��厮����V��]&�/��Y�$ г����m~��Iv����؄� n������a�\����'<#��(G�thͷ^+�1��@w��D ��_�9o���$�j���}�$֛W����%l�o����+��a¸��Q�C��y3�p0iCB*1S ���@ɣ��!��.�h�To��x��5b��b�f+ރ���8�o�˳+���!b�u��Tm��dEl�Ƙ4����H5(M%z���e���`��VL>�
K����f�9��J��y2�����1��)=��H>�,���u��۝q@f8��!Z������{\�����$�Y��Ŷ1���4�%kI�p:���B&*\��<����V�����e5H ��$�.��X$ �@�uA=|/4#H�� �"��4
!^؇�	�fn�v�����חNѰ�4�$#�7�7%Y1�@���ޙ'��@�A
λ%a��+���Nz\�K8uZ�
1�ݣq:L��m6O[���Nê
��RV>1�Im��P<�����AKA+-�E:��^�.a�-��W:C=���m���@tH����ez��L�<���6ᰳUl#�f�)� ��y���e��ٮM��5��9�#� ��rE8P���
�