BZh91AY&SY���& �_�Px����߰����PY�n�F:f4fk�BIj`���4�i�$6�i��i� ��M0�(��=LM@�F�b0 ��H��Ѡ�   44d���`F�b0L�`�D�j=D�D�G��  Ho���bE�D�4I�������|p��`�# �Q�!���㰄m"lm�A�M�mw���M�	n�۷2,��eۨpߞ�c���-��c`�-N�;U]����c���+�V֬P��]X�#�n�P�n:�Z��+�zM�$�%)DB��6K��<��0$���g�ޣf�/��i�Ԡ�`�l_N��eM���a>	$y����A���mQ�3�Z�.��Z�|��ݍ�VՒl|�	�����Ga�*^�ԙ�j��J�1�R��\��%(��#�X�W��بG�)K��QĐK(i����7E{�Z�(��.��&����4��d��vz����F�$	~��m�BP�coMW���N��mz�&L��X�&'#6;(��2@cq4[�h5� �}�Maߴ3�-Xe0ѫ�CW&a%E)l���23O?G����j������<<��?=�l��VQ�=���)�{2�%�]޾>$��BLO8��@�����?��;�:ZJ^����6��%lŨK�p�ð;(�!� ��Xmhl� ��/�H��3xh�X�D�oNx�n[M���t%��/�Y���`%7lfb�F�S'KҘ3�"[����P�Qs�^�k�˸KK)��9�صӚn�����uv�{=���tZ)��`�)�4�v��.�[ L�F�â�D�" ����4&caN�ڃ�����ނ�w�j����V��xk�D>Q!����L�T��d��'�ONa�d!�=,��b�ňh,;��6@��7�Ӕ�9 JWp���(�G�\�F��y[_[5\�Ņ�HG0%�ҷ����Zx�"��{� �pdT�ﲊ��cE�!�Rz��"	���|��4T�{b8n��Z+,�uY�(JV�p<�!�	Epu�/�A5��$FK(%�Y2l�J��F�����'&�bOAC69���p��&H�9�G�ZT�$�h#�2.ݴ4���L�)�К�g6��$��X�j�\�L�î�q	 ���S��<�;k4�I>�h[��y��d1��u��U��I�,��@J�	O5'��b�(Ё��&��������B�ȅ �n*H���ȡ����P�����EV�ԦQr8�����%x�=ƕ*2��ql�3i�w�!��-���"�(H^M{� 