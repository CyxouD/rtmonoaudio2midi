BZh91AY&SY�4 �߀Px����߰����`z�s�׼�
�$�3F�(ލI�	���SL��mFCM�5= )( G�  h  L��  �     	OQ)�M$�h4i�� �Ѡ���d9�14L�2da0M4����$HM	���@$�6� d0���=�@H�� @ W�H�C�8͏<7G&d�0� bP��N?���/"�6�&�(�ָoZ�t_�f��=���$��m�mm�'�UɻDXaD�D�n�5QQUQ���6f�]b�b�	��[H���ӦJ������h��H0E�D�+e�I$�֐�7�����3&���M���y�����cE�Z���*��	�N��S��w���=o8����U�.[6M�I4dA�:{u��q�Z̬ؾ៾d	cA2a��J&"��$)H��ƅMI�Yղ�Ԗ�^͵gY���R���[4D��k�HS����.V���n�5�B�m�D]=u�E��+IN�h �j-^�N�	9iYBe@R
� T�	.L�Di��i�W���D��B�2gyDU@�0�I/AR��(�"�a8Reu.c�D[�0j'U�V8�Y"d]�Q�,؞6�׆ n�K7�t�w
�`̈�b�Ze������:2r�Y�8�W���o�o*(��U���vy\aI˞�K׍[�0+�F��}����2$F�b�6�A4�R��1�,@!����<��s½�SZ���a�I�1Sc����g����Y��[g7w[��|	p���
3~8o���֌o!a-Tr����
�w�I[A}���B�}K;�~^�$:`a%�����m3�n#R����8�����hb��"7��O��7Rӊ(�=��L��]�mQ�#j�lћ���j7 ��Ը1���b-d���zF+������Ir��(�;]S��Ъ�R��+-3��n���ό�hA��&I�h�AF�$9���� �/Giq́B�"H9f,يf7�1\��1���R$��^Y}��5�y�qM룕A�C��}I�"RNNg���Fr)�/ͭ��l����zWVD۵��9�^�q�ٴ5s̔�����M��K��?�@��D�㾗��Ό��l \�q�8w� 2�l}���0�}�芐�j�M�P���ƊȌ��a+��D	�|+�!�V�' ό%�D��j���*ĉ��A+I��W�@�T��T��ƌ�e@#>�tsd,4BZq���2�N��4� ��Qv\:Â��5�Cy�ҕdƀC�Z�2N���@";�:���n���_�Vf\�`�)���GN�	�"`�Y����x�J��vAO��A!�j��L9b�7g{*�E� �3�d8�r���A�s,X�ۂ�3c��"�I@��&�fېUKG1�ku,�Wy5ju"�K�pv�@���lT�-��7I�|BF�G>�_���"�(HB� 