BZh91AY&SYT��� J߀Px����߰����`_-�UW*@�*I4�M���M=M��=&���&FG�EO�&&��      �A�ɓ&F�L�LLD��A�=O(  ���A�ɓ&F�L�LDI��jjzOM 5OoR��4h�$�r�"�H��% �/"��������,��G��P���H�|h���ch�a"�/k�R��Ŏ�.+�@�����=N��{l/�w��K�)�܆w"a�)6ل
"�'-��jT�P@��pH���|�$0E��
����a*����� ���I	h
C�m{�=0L�00z_��z��������X#����Vñ�� ����^��jI�A#Ŧ�J���#4u��C�q���  ��9�;�pt�zȩvv��U�
u�W��Vk%Pܰ���A�E�<42KU��pT���`QoLf�u$�Z�3����b�VL����,��fU&f��	0/9rN�C�I
�&j��d;��刁b�{��0�0�Ζ9#+
hX)M�T��v8	L��/`��5ҝ�P�^L������L��MƄd�X�ˊ�VܬjY:�s�����רi��`��-����ƚ� �  !M|���R�xv\�R�ZvDY���&mR��h��Hq	@ѹ����P~p(s���/&,��tv�&A������I3	R�,T�}�	���1�ł���~�͸%�ћ��.y�/��b�];>��)��jt( A��>��HلB
EątJM�a���^H3�)�h�C���bA0+�U�6N̷�E�(�Chp������|��^h�W���B��i�9��AϞ�<w���,�Xn@�~��X�f�g�5G<�]�)[���H�-l�{�n#�+裻+Zg ������-Mt��u�ML��P�	mbS$v� Ӻ��ƐS�
��w��E�J�:
��3<}k��cj{��5�I�B�J.�z��y<%�>=�!ʀ�%mT�U�U��
~w��,T���L$����,n �|��+g�s�1�]�[�K�?�0~w8{;���&thY�`z� Hg2��p�6vX���(��ȱ"�	�cEd�%�7�!-Ǆ���q"�2�*S�g�#���Q;D\���U�7e� �pGW��=���Ɓ�:| ���3:������?Ф:�j�vT�*.s�%گ��A�=����;�sb��h=�:Ў��p.ΰ�j��I����*�o*C�
���Ióਕ���5���Ip>��0U��ҩ�{�AI#�
��wa� ���>]P ��Av���1WJa�%R�GB�<�_�jن/���$,�ID���pU-IL2��g ��fb{F;�����Kh����2���Yl�H�i�te���ܑN$$��@