BZh91AY&SY?*'4 ߀Px����߰����`�z�1� �Ul2
��&��@F�&=2��@�4��bO 
R�i�	��� ���h� �@ �A�h  $�SBQ� @   M`LM&L�LM2100	!�)�S�j����zOP4��z�����-�$��4�!BBA�@���+�{���9�h��0���z?9�1"�m�!�Y���b�U ����\G����44!��`���;ծ ��* a��M4P8I��U	�Fh�P A� ��
��B�e��J`��Q�B�j�A�,�$#�jYaz8Xa�b��K#T��=�3�\��*�L�����b��?����a���ݾdp�o_��ǒ�����O�Kֱ�*�u��G��!�즒eFYqhS�q�}��˝�_w�M�����k�ȸɚ�=�
�3���b��[��������<����a��f�3�V�������W�S?.w_�;c���!�ڢ-Md��'�8�K�.S$����Y�l/�ɰ�L�2�v��8ڂ��K�����M�_uJ�yaJ�2:� ��,�&3�u|�N���#[jz؋B��ĝ!�����.@����Qx���L�6Q'�q�^�jĄ��6b�VCڗ�
��DИ�t$P�����s�8"4ʊk�;6�Ԓ勉1L�D,,�ŗ3T>X�4c ��e��D4�""��m6nY�]��Bu	W��]�)�T��:*.�r���xvg��sQWj�?Bz)t�;;q�I��
�a���e�})�5�{dƅΰ��{�&���:L7i\�\�a���e>�U=<N_<�������7"[����^1�*(�AUP`@(������.ON�L�}���ӂ�\��Hj��hP2q4 �)���BL3��Cd�TCr�@]�3��8��X0�av��Z�+Ci 
X��k�]�<{	�)tc�fs�s���k���yO������p�b�K
~���ؕk��N���=�䬹���WD��7i�ƅ%/Y��+>��9[1��qsh��?�~�.�\7�6̄��MQ��4mWڈ%G�9��r�7`G�`�їR����>����K�͹�3CQTsI#.�m��i���@d=���L�u��d�F/}T����ӝw�T��sו	$�Z[Q!%Q�Nt��g��P�̎�1��Pb) ,�viLӁn�J���6WH�oI�\pUS^}� 0)��7�">�"+M�W@4	�@u�x#���u����O��$�3���01�e����b��Y�R�8@)��0�\��x����Ӳ���Z]R��#$��@w���4�9���r�L1@:"�=D�z*�4ƋH���RX4!	�x�"B&(]I8yB7Q#]M;DQJҚ�$J�$�7e�* @B��K���ά��� �Pzr�,�f�T˫�zC�sV�bUEAL�9͖��F`�T2E㑸�u�J2c �q�t�I��zH=� !S쬪xe�g����LV���!F2`A�qn)0��y������>��<f�}�bW�c:�ʜ��7a��
�&M�x,��!J�2�,�_ կ^�/rA`!.ri��;.<�k^�b���d���٘�Z����q�3��h���,����ɳ�$����Hݜ�U�/���)��Q9�