BZh91AY&SY��E �߀Px����߰����`�_x �! ��I!���<ѡ4i0�ф4�2S�@M��FF #��`LM&L�LM2100	Md� =@H h  hj��!��=#&�� ��d4 �&�FS���56��=5 ��M�����*9AK�P��Z{�������Y7�p$��j�1���苡2��������'��U�^�G��R��*�W;T*&�rQ����c��ߔ��(h$"�^���i��� B�/E�i�l��؆��z�"&yidD6����wU0fdF zo��#9~�w�%�n
�5i���<uW$v�^ے����q&��\M[DJtШ9�n�,5���� ���-��)v��2��D���Z�a�]*�c|�&,D�Q�T7��<PK��ج�����R��OZJ�CI�oYI��;���M`�eMfi=��P�2[)���\>�rm�ö�6�4Z�ی�les,���XVLSN\��4ˠ�M�N��$�e�L�:�d��`�b��P�S`0ER���v�XLHg7.�kV�R��ꎢꅅK�J���3I����XK��ӗuM�5N�J�i�Q�a�jE�`����𖡄��Ô���S���';
'����X�n�j�)�n��ƤC�̦y�eI�*�]���BBK�$�@�a�r'è�|�n�;�5%Tm����z�G(ౠ��u�"`���U��%V��z ����y�:�f@�w����2J�
�����ҏQ(�O�.;5�k�;����,��*�����Fo���}(��,*�$�.�Z|���l�*R��* O�97&��D�ƚ������,�L� C���m�����=��<�$T�J[9�՜M���A)t��9?��GM[��_ጸ <�$
=�x���2tQ��&�'�>�*3=�,��#9�R�wq��B�YL\{�h��{�4e�}��ވ�@* �AG�+k�f1�Ɨ��(�&4N�Y��`�"�Pe�sna�Y����x	���g݊�'���ܛ�õPu������՗7O+ ���k�P�5O�O���0�^C�I�d��.\�`R\B91��&�� >����ax�5W0�0��:O���[_�Ӎ5vçc��Y�jXy��{ �I㇣3�t�R\4'�&2��ˎ�8-�HB&v+qvd[\Zî�>�{�	p!��fPC�I�Sw9Xs�4Udա�3{̀�^~���.�Ğ5@���j�"�n��U�0z|=%Ps�����T�k�٭��3�wS�2C�f�V0�$�����҇��7��Tq���O�ϟn�/N4x�`ujx����^^M��p���<��ih$�U���#-
���z�V�[ ������*��8��K����t,�2�"\�YeR�-�E-x�HxE'�	�5���Z�Bպ�r;l���J�"�L0pv@,C2;K��b^g{1��H�ɒ4��?�w$S�	�tP0