BZh91AY&SY��� _�Px����߰����`���z� ^*�T%(DCA4��*���cMA�(��jS��U  4     ��E ��     S�%4T    12   ���a2dɑ��4�# C �D�B&4�M�M=�5=LЇ�hѧ��*����@N�DR@��	�$��y ����~7UfXP��͔�
	4f6���,��X����d�v�$�q�-fgiOŠ�ApqYAS�8%I��0*�)�)��,&�D!����`�a���p�Xa��Q�c��d���U	��͎>��H��p5���J)x�A�xJBJ�!#!{4�u|�&���}6zU��׊������M�ʃŃ1[Hw�wӢr7�`�(M,��(W�J���!��z��`N��Q̀U��J9 �vn�U�DT�i�^A �QeFV�8�����p���Q� �=6�Jc�#�=t*RiD�\���CQ�n��g�Ք�∤P� *��jAlb,=�D(
@F�]J atNjꯜ�9��b�X�U\T�׶���Q�x�[%��y��"�l�6f�uo8���k]��.�X�[ۂ�Bq�Nz&bOH�r�&&;��]Wb�� �i�ѭnx�d��*򷆎��=Dsc�7B���g�3��Q�ˉ(�b�[�8�s1��sD�	"<�!L	r n=#u8��&��'y��ssF���	&�Y�횦()VG%눘/-��_I�.�k��r�K�����p掤
��Xe����|8&V����$݉�S���Zo��XF��	*��lU��ڎ^�(*<s�<�;���1+���Vy97zE������� ��@Aۓ�Oq){��5W�g�"̖p��P�2�G�1R� ���BS���	`���� r�Zb,���M0z�󅥅��j�����B�����D����;-�}������Nq,��z������rӅ�7@��Yӕ{  <�����%yo�b���9ɺo�o���VW�\N���##1�����W�0��.�b��B�p�	�;[՚�E)|��γ�gt��j-߫j��i�凼����H�f�Y�^aJ�ݞ��0A�y/�3;���J)�YE�*�g2r�+Q�2po��Mx��H-��#HDA��iҺ$ʐSt]��=%F"�'"���5b_�Ը��j���X�޳Am�*/���o`lև��ϣ遐 !�"!�MJ1�B�F������H �z��6����)��yc���O���_����`r���=���07��o	��F1�bc,��a��B� ;y��#k3��~�0�C���'��0��>a�4^H��U;��Є&���Y"(*b�8w�7U#`����*�A6Q,�w]��U��pO�Ѥ؎0�@n�P����G|k�0}��iV��z�
ٮwmWwb3%{$fN=���ۖ�#�L�߸6�z-6=�B�����F��W%`r�[5��10>7�#0<A�����Q�ic&
�J��D��L�+S�b�m�Mu!r��F9�[��ŀ��r裗��
n9�h��m�T��)���)
 p�E"{�p�ŷy�ܼ�gA�}��-RT�4�k���(dy�T�1/��A��&H���*��ܑN$)���