BZh91AY&SY���m �_�px����߰����`�}�}� ϗ��AI�ajc%<����6��@=@4�5<�*(�� 4f��i� M2Q@ @    S�C@�!��d0��  �R��mA�@��d 2dbb� �$D&�bjm�OI�P��� چ@ Hu�u�Fx� $�+� �&G�P~��Pe� �����	G��BYf6�l!�U�z�.>ܴITU�B#�� (��Yg��M���\�TRmH- �Kpm&J)B%CFT�d)i��RHi�
RCi�����U���VI:�BFT�F8��,q�Fd��ב���og�D!�r� �_Fa�o#���4�&A%����U���ajG���+�Q >@^PX�d�,�n�����R�s!�Gg�۪�=L��i��1��:} O,%�&l�Y��k;���Τ!=��ɠ�&i�b�!��es���Ht��@`�4�a���=f0�".<��
������8׆S�OS|Z�"�^kKC^F:2b6�d���r僳���N��N襥����r/]���ػH���40k�:&�>�:�&��o������,"B,�R�ʐN`U���b�t#��/�͙�3![�*���c���iU��Z�3��c�J�"�1eX���e�:�nձ�ΝQ��� ���šf.��]T=V ��F�I��"�닙9uA���݌�m������<$�H$�$�I �89"B�v�- �9y�*-t�L�B"��Pr- ���A���@šh�J���I�$�4����N��!h���ȷ>	!�,�b����2���h�ϟ.>Cܺ#��ɖ����'��]���9��+CN�ZT�@������(�`L�&I���W���~j�:�g+~^GQ��x$;N�z6����h4���H�A�� g,7��9O"� ����\��aGM��j_��P�I�j\���V�Ӣ��M�OM���&�4������ĥ��F/~%T��M~��� ݸ�s<�PЋ�$�[IL���N��L�;��wE�G���v+%$	΅���mĿ�m]*F2�����d[,U��rIį5��(�����Ҙ0�T��:���|�|�t�s��L��⤐.�+o(-!�y1x�m�5���H�lf�$
jma�a����:A�T��Ǿ�a͜3Z�buL		3�$Ǌ�����s���@�}�ꋐ�y�U'slcE�J'bq`��\�2���q"(.d�8}��ڤf,�U^%A&�%�N�İ*�wx\�z�:ҒzH�b(9��1�p�d����*C�F��=,�9�u�u���������iE�2H]F�#ra��m��Ir��w�u�誂�ڦ�mK0�0T���PF�6e*@oC��:鶸o0a�^Tᾢ�̜-m�m=������I���!ǟ���U.A�t,�֙b3⡴���Rpk �=Ch�/%Rװ�l,]�3�j��z�T����pv�*�dw��b_L�=���$\ɒ<�;����.�p�!ם��