BZh91AY&SYk��( �_�Px����߰����P�q�S����)XI �5LOSLG��M���	���dɓ#	�i�F& ���MI  �@   ���������@�4   d H��LS4�ɴ�F�i�CL@ �sEc��H���Q*!c�����|(���O�@P=���b��V@% �L0�)f[���� ���y��~�DG,�e�v� ��Ѝ��$CP!�. ����a�Q��@��I���0ENȂ�e[ZA�+p#�#�T�{���3�N�HI]<$$y��s���+&M�����������̻]��B�L�����])�a{�c�pg~C��m�Klk�� �o)�6�Yk�s�CU�����yţm���;Z��b
�8X�ATM%y�l5��ƎDce} ���7�mPj��*-Wj�^�U0�!UP���.ѰA��$f�M"�3�CM�@�4�^KL'3���<cSW��b�R��gZ"�1�d�EZpQ�RI�"$n��/�nԷn[�p��F0Z�,��2�5j�8��^�>/0�$��ޖ�m�@�J�����]]|�U�%�s��y#�������&֋2B�h�A&|PЛ����$��<���P�aQ����ɚ��6`�^^��z�V��p��R���}�_	����כ�t�����_]9^B�w��K��~=�����I��[L
;h#ǳ���F�����MGגe�Ƥ	fW����M�1˘S�� /�$"$�q�[0F��ZMl�d�I��$x���iּ�0�@x��R�K��V�N��":D����Ԑ�e�k�;9���S�w���cm�kâα��F���y3�poBRjM��Q�4�9�4���Ap:^�C1�ġH r����3>b��u��q����&����Fn< -���~��D|Xн��BUL��z�Bh�F�F��F�yi����`�y�bTf!9�[@lހ�Ia�7@�y�fl�m��874G>��1�|�k�\��� 7�Kv��xF���|.P����������ܮ'��-"3�N��h@@��et0B�I�3��D�²���*Ĕ0�W(�6�W��@�*p������@K|�m$�Ս��W�!��[�b��I��vd�3^�6��v��6��.H�zq��`y7�WĘ{8\<�P	9G���t��eF�5ƥ�,]��c&��N�0oոn�E-��
���� ���*J�Ί,R[!���~�Z�� �l~��R�E�9>C�F�B���He��� �Pɤ]������B��L۞K��5ۉE�JnFqpu�V��0Q��S��IM8aK�幚���"�(H5�b� 