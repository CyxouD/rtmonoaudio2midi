BZh91AY&SY ��& �_�py����߰����`^|﷧�:����c�8IDқ�Ҙ�ɧ��4����4�	4�b �M�4��  �&M4�dd�т0�F� Jh�F�@��  ɠhz�DI�)�O�4�2���4bb4��d�PH� �Jm22I�d�Si= ��=OSC�<��BT� ćg�G=��t?�S�?N��!�R`_�$�yM	,�*��w0�%V5����3�G		���M@���B�ӛt��]g��5ZRD��	�nݺ�zzFZdKW ƌ�id����s�����렐�ō$'�;V��!�� ���j��5��_�%�*�rH �q��(
��yD���~LYMz`$1�07>�e�����%��˗��3$���{ܹc})�em��] ���F]2�{!�|.��W��3D&��`~A�� g+�0ʺ3���T�ڞ�ѓ�im)-)��0n����2�1�h *����ZX��>��KJG��gu#�\����0�֎�1*h����0�%�4��<��,�2J�ѳ�� ��Pnָu�grr7|�D�jӀy�Mb��B
��IMIqQW���J�;�����$$$��&I L3A;m���$������:�T�*"̓���*��(��I�vu���:	c$0�@��iE�!���Df��p[<,,�\�O�d�1�$bы3<�1�u�˭��z�t`�3�Xs��C�?ΧI��.����������KtO��ӿ���0ѨI������*S��}	Ě$U.B3�3T/���$P+8�mؕt�s��`j�h��G�Ci�����=O��Ԗ��J���D���:�2'];V��7=��`$[�s199��QT�@S�RO��*�*�\����D1'c3*�k�k�;�e(��95��v'�?�d���I�ax�" �&��Η��{	�
E��-�Ӡ�1j@�䳕�ԙ���+7��p��M�0U��UMyvE�]��p�"9�^}i�Б).u!\��b�說�/5n=�P}z�ܒIZ���
)$-�r�H�;-��N"��[fT�m"���ǔ�����B%���+����E=J�[(${N�ڑ���S[���'D�CIhȘ�~{+����O��E�hB�+>���5�-���S5��#V-3r�ԫ$�	)��0y����"����V5�q����
f�,��M�\N��Fp�|�aO7q6�A�(1�Z˙wnR��q���s�b�l`����$��=�=��
�wJ�̶�׳��R!�\,�B�e ����F�
��a�s�b�Fz5��b�-�
ƁKe̦�E��`Xĩ�~����{��Z�E*��V�d�R��H�Ue�{�Fm�������X�bU�>L�쾿cWN������sK)m$��e[̹d>�E4H���u��ӧ���ȹ!�sc	ܼR���"�(H X� 