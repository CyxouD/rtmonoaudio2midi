BZh91AY&SY+*3 Z_�Px����������P>9n��Y�$��CE26�����4Q�2m 4444��EA��A�4�i�bhd d���J'�2F���bh4��`�1 �&	�!��L��QSDĘ�ڛMFi�@hmL�("�3��B%D�@� �u�'�Q���X��(�0���$6T 1h"��-�ɠ���ŐQ�Ř�:ȅ���]7�Q���ۂ� �6��M��M�:��h#���W�8W�<�)�/&J� ��/��݇USi5�6��:�� Q3&M���^8�;���A���E�-K׭�ٓ���68!�����Va��gP�r�Ș�rh����1���A͘�S%9��*VJ1�U!��f�,�!��b�b��H�Q3�j�"��D�h8�Z�� DBar�e8�/JC�f
@�`�j�,�9��e1,"".,a2�4ع��@�������q�,d��!�(�VY�*6rt0<韑�i-�(�U"�R��٤itp�Lu{�z=&��������N��y�\�%�DQ��DE�Oe�jm2�00LkKAO���g���5��5����X5_2��!&d%w��ۧ��e�]~{��:='��vj1�y���O���1a�Tu�}����HH\'�w»��B��㇗u��W�tG�	J���zO��{� %ư�]�n�t���'�v��k�r�)��*���R�weɨ�;	��ÿ�� ����(��V2Í�E��Q����r���g;~�R�;�db���ڍ�&���a��.���n�F��" �"��2���F���h����������Ƹ� �����FC	l;e����u:3�Un��` Q�x�:ۆٛf���ot^�l�.�F���e,��Z����r]	�!B���Ai��Rf�u����'$�L qGY�9�,���HjH�g|���v©j���?��P*X���/�cq5�7&��VJZi�)p��P���5�ff�$+ą�R-<D��mk�w�#Py���[�_�ƍ����Qdn6�M�a!7%��6&�Z�W�	������͆��Q�*�&�!ð�D�A9�:0/���b��U
��	��K�Vj�C�Lj���HP�t^�}j��(�h�)WW)k��;<���`��odX��g�ML�i��T�NE�8�ub��ˁz�~�u�y\�L�T���c<���H�
%eF`