BZh91AY&SY�}D t߀Px����߰����P^�`Î��t�k��H)�6����aF�H�j=L��4��jy��S�h)�z �   ���1Dz&���4 ��9�&& &#4���d�#�#S���OTx��yM�� 4�44� �ߕ &Ċ�BII�����?o�	�6R˰l`I�a�����ch��El(��Kg�/[d���I�t���CLJ営�S��a�� �����d9����T$f�oo1��`����y�`����Pfx�I$^��!B��'ô妉�M����3f�yu���������`p_v��.��@RHB��<�*�"�Di� m!+V�v�0�&��o�e�J��&�Y��_/�P�S���¬*���U�L����h�A�Et`2����J���N��:!қ�W�kL�$k��5���1�mj�����lm���v�m�BPA6�������UzV{�d��"�-�`�H�V0�k�\0��a0��2T������]�����o��A��f���eGTSON[p�;����[軖2~�7�7w��p���;m�W���\�����N��&)�}W�^�Gv�߾#ƌɽsS��twH��̄�+tU�7��@�!pE�C`�"7����c�ןj�Љ������m�����4W��K�1�H���)rK���0��N��H�q=m���3r�%���s�Z�˓U��|[V�Q���v�;���3�~=N�2.1M%2Gp	�k�Mt���,���`q�T��Iβ�m4����y�f1���I7�XN˪j��x%t��kɕA�u���4%)(P������SÌ*V����d�n�����V�"\1SV���WF['|�U����;d�� ��D����ogO2�;�����_��Է�l#��nz���T\���aDj��;��y#|�v'�&��}	@U�Jp脻UH�Z��UM愹&B	��g���*�rm�&���X�A,����:3�a6B{"]^R�o����'��5�sg��H��$c��۩*��K4�5�I��A��m���W��a��Ͳ4�R�n��"�õ��B �5G��6�V� gmj���|h2�uZ��}��	90�����V΍Ѿ�ѐ������sR�\����� �����;@�W���P�u��A����*����\���	`��ʫ��}|Y$ٮ!##M#=�7��ܑN$7�A� 