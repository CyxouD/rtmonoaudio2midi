BZh91AY&SYA�V� �߀Px����߰����`^��׀b�*��$��$��Bbhѡ�bCLL�S���F�     )꟪  Q� �d� �	���dɓ#	�i�F& ��T�  h�   �  ���I�S$�?MS�zf�����Hhi�zBg���xO� O  `$� �1��� G����U��l`5,|YH��PI#�,���a"�/k��l��� ���T��5`b�8
�CC)HAnBn%Ȓ_=px���'�H�v�&8�,q�F<�3-&8��_=�3}�R�$��[j����:�����Ƭٺh��n�{�f���k����l�{���	w]��)�,a18V���2��1Z�$U�,\,�5�$.�p��x��{R��,g�
)������U *iE�l��$(�И?�2!iE��RPd��.fkaN�۶�8�.ōF�*��Y��]"�Bƀ��dqHV��ډQ�eK�n�ԹU3���P8��]�5�kF��0�,�E�2-��#X+�����x��b-*�Ôy�|L|�J4ذ�C,J3)y�٤g,���M&�6�ĺ�Q!�9W�aI5{S%q_�L"�(m�`�ϳ��۾�Ъƴ�����[��N�4�v� ��t�����:�cco[m���n�R�R��骺���d��"�E�~�`�a
A�"a�v1*5�h!��CQ !����P{����Ʌ�Wxi�H�W[�k��.�r��\{��9��]�nBy{�W����9?>�-5����ZW���`���G�w���j�[L�D�f�-���޳��8O��9msPԵl��8\�P��]�>����Bܸ��M��b�J}*/�NX6sG��%n�����<�I��.Լ�`�02tQ��� ������=�v��S9�v�N	�JO}!d�L�sKMZ�;vSK<�G3�-
� ��H4�[�ƐSl�n$u�ʕ� �}�o�1u$�,\�-bU�P�k���J���� "����23��Ύ=��K� ��ȡZ7�z������/(��J�	����C���W���fo�7tP����k�����61间����N:��ٱ�&h���4�G88v��4B5��Nױ�"�����.D4	E�T'�i��3(����$@��+�$E eKԧ θG�T�z�wDU]��e�Gr�X@"�	پ�O��#J9 ���$Y���^�ן�u�<�=Ĭ�Pdi�~�;�é`�5��Iá+����HD�'gV�\�TqE�6���F^�^{q.D��4�c(5dV�*�=��x��o�x�����V6w�k��`�N�3|� # �e�*C�\UQ�����B*�k�!�55�1� �$#`���X�� b�꩜#>�p))��2�pvA ���cTI���d{1��##&Hޱ�0�_�w$S�	�k�