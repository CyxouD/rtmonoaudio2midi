BZh91AY&SY��� �߀Px����߰����`�S�a���)
���H�4����&&M4��z���jzA��� MI@�@  @ �	���dɓ#	�i�F& ��#R�@����D  �	���dɓ#	�i�F& �""h��A��CJx�&�Q��� �� H�	1"�@�I$@�p7[�!�~eQ�30"PB9�C͊D�A �sG�i0�������F@�sJ�t���
:n"��謮�8��+X�b@٪��7D(\ � �e:)C:�O�;��{@��*��*��	vg��_M�ٺx��~�I*R R/|�M3�i��32oL��Ça�شv;�}N��87���~ m�]�M�	F��B�[n���K�K�}�y*�Е�J`�=V"OM�ouJ�l�4�i"����
���#69TI	�k���� �0;�&��QyR�֪e�T'&Ȍ���X��m����U�`�S�O҅mx�ft�ݓ�913�7$v���%ʍ4�����ֺݱ�;nl���D��LT[�L���@�@�rD&��4Z�����i˖����1N6*egr�,�^���4e�8�Z�d��jI�E]�b@��Q��4��Jem/X�,t�Ch�U:ޘ��bg3]lrl!6�l���Wf��ɻ�w	 �I�I$B�w�m��:�?G~Չg�J�28R�����G��jJ4Ht+���j�A�%�E��1|�*c���(X��a3'�U��3	��w{��i4�Q�z�]g��)���>є�o����?~[�*3��=qm���pB<me��w����b������A��r��C>"X�v����ɳr�U��ˤ;������xu46G!����Rhh�hVT�����(��r��M3#�s�-���1����A�엓xj妢��JEw�WӜ�A0�޾G����Qۍ�3����]���yf�j��魞����70%�xĒ�#�:�	4�
vAp:�G�`tbTiU�!Β횓5`[�Թ=�5d����&kE�N�Q�=��N?:ǁos>�+��B2��vK�mS�:nخٸ(>�r�W��v��]������Θ����1��C�d]J�o[�f���͍�z����0?*�8{x�E�,��fr�M�  B=�Wz�������}Na#�TX�����/��<�Lh����U;���5?�$E eL� �HG]R0��*�Q�2M�%����\!rx;6�A6-4���B/��Q*�ʅh���ä��~.�D�չ�~��c0hV2G1�8�����h�B8�K�vu�`����Rǟ�_�-&��Wi\�b�*k�P#�6%*@o#��o�u���4�좵�*&�4�}�b���U��,P��Oe���vD�=�-H��Sb�B�V��{0���}䅀��(�v#۬��uq(r�Z��8AӖ�압������zQF#h��l��.M���!#sM#.�(���"�(H�e 