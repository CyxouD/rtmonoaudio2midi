BZh91AY&SYe�
 z_�Px����߰����`Ϟ%�c�"�%$	$��h�hЍ52h��	�i���d����A� �44��14�C@sbh0�2d��`�i���!�i�MA���z�    h�	���dɓ#	�i�F& �" �4Q���S�=)榓ڠ��OQ����	
f �9JH�$�'�|��_��eF]�`�! MC��Dƀ��"�mXCH���]��HM~��(��JI��)t��}k���ׄ�k�2��A.�&I�P�Ba!��dd3 � (��eb����cJ�*+,c�'`��h ̥ai���Ww(�W9 �\�����V	�lyt9n�࿭n�������7�����`@�DM"(���@���4�\�w8N�p%2>�%is�=G)�;P�U��D;M�z �!���Pw�ˡkK'��!m��9���[��p3���KF����/S��g0l�aq�]"A�|�¥��[�6�"S�0��a�
p�.����C�P�r��=&�֭�t/\Hy�*�&@K8�1r8��T��`�MB$���%5����v��5���s-qO%���V��R��jӾJ\kmL7"26Y^�3��
ׄ'Y�U��)3�!X���]��O�(}
ك�0n���_*�>��N�]�bCDkv����'��6.Y�Q0���\WRz=|��  $32M���z)}��j�R�jt�]��˓7��1clen �DcX���X6�����L�ā4��*�����T,�\a�Q�����Hf@T�LV����S󒞚y7�Y��\s�~p℮�W���t����1���F'�V���! X�����Sf$�*R��
 M�1->�b<h�T�}=G��q���D�/2�ϧ�<.���J���� ^�f��f�5f�ͭc�J\�g��7,�H����i�z�of@zˤH��x�� �,d�ѝ��O[9��"�oIu�h������{�8m5v_Yzy�Ij��Sc?@Ј`CBW��&H�A�Z�&T�� �:䎳㤨ҫR$	΂�sL���k��c=]�s�6�jhS(��A0��g,k�&��l�i T�����eLQ�ە�s���)߂�6Z�|r��*7Ac�D�1co��a�%���	��;�K�����"q��\���~��'�aI��@�w.�3�s3���P2�Qrd��T'X�-$j(����	@�N�U�1�H� ˙)N��#}R4D�Ux�P �(�s;�E��(Ul�� Mv��7D�\$M$�8��,4­Qm�Ҩ9�o���+-s�-����¤�����:��Ņā=�8!I��]<`=�@���g�tm'�]&��JA�Kp�0�Rp���!vx��ë9��E�+�,d�"��}k��u�qو`Ic�N�@�b@��M6�#nJ��f�T��в�=b6�����Ҁ�A"j��j^굣Q-�Y�/�1=�J�#%�l��@�3#�ȣ;��sَ9"�L�}n�)���"�(H2ҏ 