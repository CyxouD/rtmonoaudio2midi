BZh91AY&SY9�- 4߀Px����߰����`C�X($$Rhj��i�3JyOI�544��4mF����i�j���       0&&�	�&L�&	���`LM&L�LM2100���&L�20�&�db``"M4�'�~&�aG��2���hU��2
� �$I �	=���$]ԩ�&�(�0�R6(�!CGC4�XI�zV�*�H�\x\�{�y����μ�(vk��	g_�1Ir��˒i.J�Ud�nD|���3�6�JJ��-L�c����0H�3��SI���?��@V���B�������I1 �;��*��y�?c��b�_�mp�x{�=1M���7v-�s�*�+3#�|^J��7}ci�t���N�7�;XD����h�B����TE�d�E�8����3dA. �.��xa�Vq�l�MO���̘�%�\4C@Ȉ)j��gK[)���(r���%:���8�/E�D�R&;c4-�c��j��Wb��N�D�Ӊ����ф�J��E����$4��m���T3!��f�ma��eWM�}hD�(�H�5/0�H�^f�H�x����1��h;���3�:�H$�IlH �x�S���ۻ�����DY��،-xs�r�� ���kL?F�&Ҙy9Y�.$�
�����,.�I���ץ��m"�/:ݽ��?T�WFL6k>Ke'_~1�m�-����6���xv�`6^�qa�累UZ���f�ߒ�0��c���(�n��g'��{�閊��_�"�g���,�m�p� �Q ��� 8@�?P�g+�ʱ؈�.�D�#�
�ÚH��ʨ�K�+�3,�2��j^�X�_j#�2D�
d����"v�k�K��6��T5WM�q��4���~i��v��{i!�\`#���H��N��L�8�`�Ў�#��Tb+"@D�[�Zf�K��7�#P�}�Ħ���eE�����r7Ͼ�E���LH	��Ht*`�6ڭ��(>�r�8�1d��ѓr�61�b�Ngc2&��D�`�-�Xt�@Wf61���y����]r�ś�-P��F� <�~���F�ٙ�|\�(��:��4bQz*�cE��e�84�&��}$����Jp�!.H�X*'x��Ĩ"��D��	 !T#��H'w-e��$A =<�(6i�X(��I�˧�W��F�|1*₲�A�n�a�I�c ��Q��+���.�#�2\�Pk�$*�m6=��t���mbY�n*����͙J�o�C�}��E6W0�ц��E|8TX�	�p�]j�;�	,o�K�q 1b@[=5a��U�
nA�t,�jц!}���}a�!p 8�H���5Z��"b���S��_T�A0�@;b��Ѹȧ����t͚���i��B����)���h