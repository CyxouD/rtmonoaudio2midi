BZh91AY&SY��EN c߀Px����������`_{��z֛�ti@�I���T�x��4�O��F�P=�=��@M��F FL����L�4h     5<��T� � @  h`LM&L�LM2100	#@��Oj!�6�T�hz�4cS	�  �&!	@$���|��} ���j��0lD�ԟ���B0"�m�!�U��u�W��N�A~4� �/� 924o�A��'5=��LX"BM.I&	�b��Έ.SY�$����}X�Z�j�8`E�cȂ�
Q���6e]�bQGi@P�BY��A�m���E	� fL����b�5���፨g8�@��	�L�����IبǕI�0�
F�]9i,)�l�`�Mca0�]��"��A�7	�0�L�,�u"9&����6��bPĽN 	i2�:T�:Kv����6)���P�1A*E�C8)���xҶ��
���>S'2�:!��K,��6M��J�&K�(�GU��,E�Pp�WQ�J�Nrct��q."�*$ ���2�e���PN��3E�k*�Ij!JC���c�R�P���X;Z5sĜ-����ŮL͘f��n�)�yA����6C���3i�b 59T�6h̴m5j�f������/A ��I$�bA���R��K���QZt�\EY&vDR�Vh-�p^��q��4�4�����M �d��\g��p[W��asT��I� )�ʚ���D��'��`诨�-s��nB|\/�~�У���~9NVS�+�5NU��5B�����J��X��H���?	��������TU���3gւ�΁6����7Y���؋����?�3:��&���z�눊V�����^�ɑ�=��χ%��̀�]�@���Y�8�b�UH�����,�,�*̗�`�8����͜B�s�4o�ȶȕ�n���τ�`��RrbW"�4�9��N	�C(�du�J*5$��ߥ3M�M+�F2�{�ēzL
�z���k@���64?����y00��p�H7)܌��Wn��y���	%͘��_�n��k�P�3�2�,�M�j��x�3lcc�6C�xlG����X�J���}�HƁgZ���������"a��A�!�ר�.��-CLh����Q;���5/}�I��z�p�B8�"�\���V�� �UQ&s;.EA!P#.�|���l@��=e�vp�h�n�׿�/���\�b���|�×��\�#i����$�&4$]R�Ҙ�8�g��P u&��o2~��l��0ZR�7-!F2`Au�'@��]�q���Zh���:���P�,��P[�ܐXq��� A{@����{�Z���bG2�F��^�߃�"����&�\����κ�͓Թ`�X�+����IÄ�13���nT�q��c��#&H�P���H�
��