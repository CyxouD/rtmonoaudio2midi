BZh91AY&SY-?�� (_�Px����߰����`��� �  N=拶��%Ih&���~Ѫ��?�4�6��&CG��M���AJ�       &1	�&�1� z	�A"&�%@h�#F��C   sbh0�2d��`�i���!�D���O�'���==)��(�� hG�w�k�(���UQt��T)E]�
г�~�_���b�@��X��"�C��H���q�r��o���7��f=����Z4rj�NjM��K���9��Չ�3�8�8Z�����u�6�u�u�Cxa/,�!{iaD�Ps���?Ή&	3�_�|8z������ۘ��v;�u��Evgz�6-��ؽ��m��SbT�>�f���͓F��&7q�QLQ����/)���C��|u�[�7vP=�%b1&�=*1�j�3M*��us�ҝ�FP5١4�l+�;ǘC�VgÎ�#ͿǒTN�&2�4�f*"����^)�hh�9R
Ww4�:]�˛�\@����@#��2<�W�����,��y1�>�=S1<�T��� �B� ��|P\zH�t�#{k��p>(F���<JB��lX���˻�b"��SM�������������F��Y!r���w*��Ç�#�[�sg�Z�#k�Xm��Y��M��3�c���#�a�\8��t c P[ږL�B����,c��Q�❝��,�4'C��}�5���˧#�'GP�Y;�u�˙��Z8���[��dgn�C�kQ�-j���_j�l]���I(��yʩ�->���.�d����7�������ˬBV���Ƕ^�U!�yAc�#8�-��۶��	cnhe�ҷf2��C�O�A=zJQ��O��3��^����G��o*���=�I��<�귰kB��	��y��$(���y�����^��DR�� b��J�w�dױ6tS6�߼��n�Ds(ގ�i�uK�쉅�U�<�z����y���m{W����Y56�>���3�y�}2��~�c����zNV�w�)��^9���'���j*5Fވ�Sg"�`�5��01�b�]lO%^Zy�7��CF����w@���E9�o�c[����o����������6�l%��e<$����{T�"4d��Te	_tU� P�T�oT�E��HQ��D!�JCu�b��1wQ�z2�N�3��	�"��a���D1o�$�����# 
\��)��>,����TAPʜ���&Y�V�@!/�ܾ����	T�.�*�5�v�xѰ����y����Dَ���)��)����s�� ��R%>�P�Ǟr�X�J^�C�C.��J?�Т��^h������-����p�&����$Q�O]^���圗�&s������^���Ȼ��50�{'"c�߄>���#�6�fE��Z,�N�kh-���To�>ܲ��� !&}�M1:�zɭ��&0�6y��k��-��J�������pr�~V+��],�-��s�P�5�%F^���#�RzYZH�-�J�� ��"q��|�>�}9�������0�=�<7�vDs���5���+)�Tx�$$�	z�h�x��C�r���hO�&	�Q��<�q/��"gb�.̋i����԰� �0�8q�6���
��)^%A
-�V��d��"���{ۘ3��y�t ��	q��Ḙ��k��xJ�����v*�m��T�ÿ� u�(�����ϣ��w�q�ԉͅ���8�-8y�'��ˍ����F�zX��ի���Iø��� s^{--���&3���
�q��,*(�R��MO�f����p��/D���dQp�(S���0ʪ�1Ґ�'�(�l�K�y�1��[9.��S5%S���8>@������Ļ���A���Hѓ$ks������)�i�&�