BZh91AY&SY�.�� �߀Px����߰����`���� R!* I"hb&����zM��2h�#M0A�~�)P� h�@2 @��@挘� ���F	� �z�&� �   ��mUh�i� @   H�2E?Si�yOi�mSO$��=M@=&�".� ���HO�� �3�>���YK.��E�Bj?6S΂BZF�Gsia��\�o&��B�J߾�����L:z)�s�yZ`��z�*R8�x�B�<(�ND��w���D(I�h�Ә���2Z!1'���wl 
f�fN5��v��P�xW�R�uu��w �*��!�tH��H�t��wy}xL&``���=��6iXf��&%hYy~n�yy�����s��#&�פ�_O�U�Q26~�a�x���(q���6�(�)vwb�0��z��cԆn����[S��@��vQ��EP� d �(2��ⰹ�q���Kt�RD�!����٣Y/�f�0���z��ޟ{1EL�dV�;|6�����V'u0$\�φq2��ĥT�l����f^�$�D��qԴ�P�ml�$t8�R�tr
�mC+V"q{��0�����s�p��$C�u���TQ��7���}�I	~��#"R��1��u��2�#0FЙg�v��M� 7E���e�;�����0j�^��b컯�涜/���P�=�}��i��M�m��n]�El��8a�ӧL2DƼ��k���[9.�n+bڕYU+�͔��a���γ@@�� !�dΠ�wt��%/�˲�����Y��1�ภhVh�����R��3� ����(�#J"e1@���T��G|�d����12@��J�T5-_v�'Y,����e�F�C���ɏ�	G�����o�Ï=����
t͕Ju�kޝ�����	��zh���!�7�|�

��I����fٹ��t���|�]��ohl/!����	�:�jXjDiC�9��r*��Q�:9kя2���y~o�R�K{�4
�:�锊��9�Ԩ0&�/���x�D�E�^�:X�g�#��U�C�r�Ɛ4�[�.X`bH�#�:Wj�������"�UiHNuۭ3^��Mk�Fce��z"Su��2�D����1
����+Ǟ.i#��02)���:�#��U��
���Հ����̄�,E2b��fA�����>�LVB��
T�0�V������7V�O.�.�1S�9�#sI	u ���]���F�g��"��|�!��J/EBv6�4ZH�Q;��%j|��"(*aJp�B7�#@����o4%�2M�K6;�aa*�u��	��RV� B�md�6g��(��F��W���L��=ns[^��`�X#�p4�:������i�_���Q��8(?�(]�)��.;�<��:�*\���D�f���B(�}�GE9+��a���+�}DփQ�Jˆ_F�7��p�0��eJ��J�5�܃1вׯV4.�_9�!p 8H���k�R�s�"�vN�Au�dw��W#F<n�H�fG��K�e�f4���d���ے���.�p�!�]y�