BZh91AY&SY�v&� �߀px����߰����`_l =�
H!(I��l��SL��2��䧑��@�S��?M �!4�4dF� �F@ч0`��`ѐ��&��O�SL���       0`��`ѐ��&��$�"e=Sj��<5=Q��4�� �S��zQSH)t
A�B�Y�>�D���-�	?�D�@����A� � &a"w@��`k?S��pۼQ8����-����_1�vl�S1�G+
'�����H^�^���t�:Ao��� ��5�#�=(s$���/(�ߨu����a!����άq�=:����i�)j���n:�|]G��o/էc(��	`fA�������(z���DĢ�4Ӵdމ�L.� 'e���7B����4
��� O0���jP1��mP9����1�̥N��/]��\�\l�ve�lP��"j���q���fj��+��2��x��șh���N��,�Z�'����'.��w��kP˒�ޟ$�v��e8��I�f(PѭUi5�m���Ƶ�rI�ÄȽ�w9UV�ڸ�O��A׭l!CV���DƮ�-�zZ�gɈ�hkWM3|�����RES%y��1K`1ƞq����,�P8 ���E�w��ye�>��:_��-UX�쉲.�R��
�Uj�4@� �^,�����%ɺ���Eu��}; h@�(�--� �a��b����	˸�������z�˿��|'���/���um���h4�<)���%�d�$"���x��W^��50��`Q�A���b<h�V��]����k1�$#R�Vpo�=/�S��T�IO/P������%�^�6�~zw�L��]���cT�}�B%֗�l��B9^��zn�6ԑ��{����JpN��)=�v����Y�=���L����Ѐ�DF�;-��kcm�U��2q6���H�CĄ3�(�BcE$���.bU���mER�P_�X��H�Y�'�o��3��Á�B!���(R�U�1�~:��acaH.�u�Vr��ĉ��̀s��-�Ln6B#^��K�q�����æ5O���W8)5�="���H*Onv�=�-Ip�N��M
�p,:]�na6+yvd��@hco7��C��A��˅6�٥V*�p��j���Q�Q)�W����y�F�!�ʢH=�^\(e
�~8��b��&��jV���sl�;r��M�5�G�v攟(�5��oZ'kJΰ��Jq�6��x��ʍ�e���桠� ��s_Y���kN�f�r&�f��xAJyDT���gb��4�&<��֠HD�HDk��v(���!ţ@�]us�4�MM���xI'd(�lt��Y����;�g �ݥ�)�h6�p| �c2?c1?���f9�䍌�#��{4�_���)���5 