BZh91AY&SY��4 T߀Px����߰����P]ޗo�7��t	$�CSєʞ��B=�y�i�j0�����M#S�H���1�0F�0�	L�P�����O$�4��� ���I�        E51G�55(<�č= � � �3T�L@�	�Bx	&�3��{H���H���B�����~h�Q���	4�0����7�0|.l5��L)Wa��X�)Պ��-:�4�.i��m��4�ϡB��QD��|�B{��"7��o�V���>2�ϼ�!"��	�\lS����`00x���f�G�R��_CI�+A�s��]��}K41q�׌�i�횝�jF�� �$��?�QF�=3J���L���e@��R�]s�G(� �NCX^�`�B�I/���Hf�P����R�h�!�efa�Rd�bfҗh���3�{z�l�Pr� �;��D3�E��{���BBKJI$�@C7����&#��ܴb�:��%��nQ�A&ĠC��!�PR�!�H)K���Ahɛ)�Щ��n�;Q0pFg[�ya��=V����.��+���{�U��y��F?�|ŧ�_�q������^���?o@����@��b={�ݱ4j*zΞ�'����q��_�f�kÔ��1��Ṑ��@����V~m�>UȊTsS>59[�8�#�=ߖ;���FH���)�����X�,d鑓�#������3�k���g;��JPN�W<�}�n����2��)���%tQ�LQ5GU@��Ҁi�x���H�����\���D �e)�����3���2�8NP���KcTW/�H>���-q�SN�T��Qb��X�Љ��M�!��!�zZ�$�^��&�W�"m����>�t�h��@�ZXfml�-@޸�}�Q�^�-ε���$@]���W��u�q$\ 抒h4*䚙w#lcE`�b��F6�Q�r\,f������f����su&��W���IL%������NDhjv�ʠ�墆p��!���;$o�v�\Vhs����birH�;�1��b��F��r�V6���d��$��c�q�^�A蒅��1�;-U�;(������#Fd�+�V�)�EAP�暋�ѧm!!��tZ� ��(�d5+���i!R�h�$ӧ wuMX�`'I��0�Ӗ��0��g �a5�u'#��� U�#��Fv%��NrF,�#*��}�W�.�p�!�a�h