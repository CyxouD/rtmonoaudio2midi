BZh91AY&SY���Z ߀Px����߰����`����� 8qN�@��I!���4510��z���14�&A�~@U�d�&�И�h hɉ�	���0 �`�0��D�MM�<�4��@P   mU ���  4   ����������SЀF�=LM%�$}tA��!~IE �Q�~��K����˰lPBMC|��T��ch��E�fk���٫ ��e[����@U��vWc��9���EƤ�\�@�\�j$\C�:@�D�"TH�	,C�aBg,� �e�'�A;��CG�>k$��=�8"�+����j�A�f����ѡZ��4QgiI	�� ���0iw�-LI��dټ}(�ރv�ϭ�MsE�Z������,X�����!A�8☕�%Q��O��~���hB%[�� �	ynD�{���a�-ߣ�7�4zu�8��kW��T0~���i�S�\����`FTY%�%�^��
��¬L���v0��8�x�d.v(��� �w��q�ixӆ5�8�`�
�B\6ӱ�Ԩ�.�$�S�p�P�MӞ��D��Bpt�r�]���>w�=g)�4G]_�
թk���;z�JC�(�U9�7)F�x�f���aǝ��Bl���D5�&aVT�'��1ND����A:�Zu��PN0�����̓V^����g!*mS�6����5R����;��>�-�~Q�a�ʊ�L�ʭ������̊��m�oh����[mb�g��>_��66���[m���	A۫j�ĥ�z�5W�g�E�,�Z��Xf- �d%ɂ��Q��b�H�F
��@�$�ͅMstw�L35_׶@�IRʖ*k;���E�_�a�n����|���)����|���t��*�Qc͓i��B]���xxW`��P>��%픓m�މ�%%/Y��a7~"^f �%}k����fm{C�J�{C`���@�/��MQ�����<��)�i���i�Ty�����r�c΀�G�!)�R�ŵ�'J��H���SU	ZٷM�+�ӆX��K��;Ey)�őY�}���g�H%B�4 >�2Gh:�3�
p���;�F��UiH!'9�u�L���%�A�c-�����b[���K�������#m�0hBS*�%�<�T�q�ـ�����I[o�Na�
��`�/�7�:��k�GXJ���Ǯ_��l�R'�������0:f ����P�����s�b> ꋐ�y��Fj����1��FE�84 .��k$E e�T� ����řQ]�T�h��&�%�.�İ�%
�9����F�BV��i2�o��ЧD�����!�&��r�����9�Y�8��+$`��Q���Q�I�S��0��x�i�ւr�l����&���|+�֖p�i�c*����B(�}���Y$n�6ƣ�4n�S����ԦZ!dBR�R��7U�	`�	[LЇX,�0ɒ�r#�e]t�p��61ш��	�6; �U.mDXX���A�}yI�ZgT=/��8:��%X̎�"�f#����Ʒ9#+&H����
?��H�
3+@