BZh91AY&SY֜IX �_�Px����߰����`^.>�|� �ϼ�V	�!$�dЙ=I�&���2FF��T��*T���ɠh�2d10�(4h�#&��� S�?H�j����M��4� D���S�?J<��~���I�i�@  ����F��=LG��� Ơ�Nm�@/�����Ag9�zW���^�� '�UcH�xV�z���/����K�a-ν�)�$�����c�Âl�)�������DK2F��e�m��%D�@�ҤQH�l�AI#����n��q�d�f�|g�C�@�%z��8Xa��33A]�y����A�,�r t�=	�[���rL�I3�>�A�]���.������$�ڴ����Xa�}���"` ��\�!��w�,f�L�vQ,1D~)J��M���6ᩁr�Ԯ9x �	�G�2�Š��a-N/�ʶ�	���{�)�}I���ں1���ގ5	,����ó;��7\E�;ME[�Ș#K���h�!܋`LC~��ț����V�m=mk��y}s2��Y��
]ݑA�f�I��&L�q	�C,����Q"@�G$�V9�K��#�P\9���!wđ�&����l�	���ƪ�w6��S�|$�H2`͇�	1�	���#͓�ٹE$"���E�6�c�۾�T��=�Ρ�5���,�q�US%-2r�6��5>�:V����\���`*U4'QP�Yh�ޢ%0Vj�
�g�:#u,��r��bY�!	l��L$m�2�i����H�ۋW�{�[�KY����o�\  @t  ��I&L�w����X-��]J�E�,䈭@��\?�0jG
2�I�BD�""�u1b�KBFqUX�p,�C�+-���0��GT�!%ST�mwk��I(�O>���v.X�~2e���W�_�<i����9���FW���$�K-�����)�( ��MP���vk��jH둔�|����y��� kum˔9m#��s�8j$�����39q�VlhplY�D�Mҧ|fr���$y�6����lځч�Um�_�7�%M1���4f/[wX򔇹oIvgg;��JPN�1{�
�Y�$�3٥*�!ۖ���H�1K%�^4$��;�H4�[�ʐS\\Q�0>ٕ+%$�s�m�)�p.�i]��4�e�z���b[��ΒI`W`p��?z����2�J'��}>�j�J�M��4��?Ņ���\�w�*3��͸��b�����H�kM�$����3�%�?���*D᷒����,���$;�$�݋�0��߸�>0�#�����Q"����cE���7�H��*�8j$E e�*S�g��T��z�wDU]Q�2M�K7]�i` U����	�q�gF�I%zI%��(9�e-5B��ϣ�U����W�9Ϳv�`ڤ��#q�m�(����<w"w](<;��5U��zձ��K~ʋ�c5*��P��Ið�Q	��Lk��t�bI���a񂌱�T�iV��������2�U�*���Ev3f.��8\�Ë�:�ڥ@]��[H�HxE'�	�6���U�u�3B�꥜�/'�EI�ѐ���  e"s�=y�!�J)�b�������ܑN$5�V 