BZh91AY&SY<��� S߀Px����������P�9n�qD�l�A$�d@�Sj��	=�OLI�H��M���=�	T� �  �C!� ��*z�A� h2    �@sbh0�2d��`�i���!�H���M5 �C=I�=M��@i�����t�bD� K�BQ�|�� ��z,Se�Q ���~����J�,ch��E\����~�%�{Gˎ*Z���ՔIސ�9�JW�d`HA���\Ð�Fh�SH����'�p��	x�bIV�Vw6��:��̤�H�]Ն�:����@&``����;N>����Hw6� ���o��������hA���-�a�!_9�c���*��� D�@��vp���I)��z�������䃬�*����KT��Wd�R�R��2�i�Ȃ��iD�[�YLM�6�u�!n���T��(4�+�I�M����)�#�,��B�� �ie�zv@�`�B�Nh��L�����*kX��$c�0�^	fA@Sr��5kG"V)a����g$���BI$��Kt�9Hf��ܛVS���D#������bB6���QQ�br�����q4b�m�酃S��(e� HZ4A�˝�S���������댏����礯���|������E�~5ey�E���M ������[� ].+���@��zv��"x�u=l�Y�93-f0+���rv�o�z��QP͡�����]|bxo�ȻڑD�ޜ��9q=�#�
-�͵z_����K����v#'P��Bz�ʄA���x�g;��JpN�R{�VOI��Y����윆���9��C����[R3�J@ӥ+#D������*p�P��9h,ש3��W2#����=3e*(��B��y $su��������������	�.T]x@n�$9L��ɂ�Ϭ��@�Y���25���e��Ѵ�@(ס�a����M ܢ9���S��5�\�0 `�]|-r4�����g�
��ZCA��4]EBY6�4["7�N�w�$�MK�v�B&(UI8s�<TH��SV��EbL��9g�]Un�����ި2��XfF��@,xAѯ9h���~\��S`u�n�v��3gs��8{�����Gq�v쵅t��
ee��0G�2N��dbB�%����沣��#Rʕa�k&P��"�c��@�9OE��vR�f��<��=�%c�E)-�ܸ,/,7��� ��
�$ɷ��b�R��H�X��E�������$��4�0̀�V-��̽�3�l�n�ST��0����3#�^�&'�ѭ��9#[&H��ܳ_���)���