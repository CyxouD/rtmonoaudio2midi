BZh91AY&SYb�B 	�߀Px����߰����`�=l� ,p��T" I!OD�ML&�@O$�zM=F�1j��i�U*da0&��& 	��C�0L@0	�h�h`ba��4�       �0L@0	�h�h`ba" ���zd�b��F���� ��4%	�ǝ$�Y�IA		�
���W��������6�P����)𠐅��ch�a"�0k����qe�\���%�� (������f�A�  _-�k1���%IA�)�,q�p��	�;����V�6�ރ0����j�"BK!t�4O���ߊ`&``���,x���hG����f�>�X�j:To��*OK�'T�4��x�� ��5c��m�B�b�b��Wu��5�f��%�U8��0r܈b3uo�"#���4�I�YYз-D��7�ڭ��Hԕ�7�`�̙�n�u�'t	H{�SWPs��#�^uQ�5,FE����f��!�/��	�z<8u��l۾�uT���t�L`
�JO8���Ñ���3$x��>ٔ@�:a���C�$�.�r��H���rp��+K ��D�h_"%��#X�_+�O$�v�8��
�"���8��5r/$2�\.98���Vm�H5���'��k]�ҵ�;V��Njr������)�ug�3��[]������o��y�j(<�G{"�`�;�u�h�2�Ux���7�+NR��Nh�����ֶ�����k3��/omP��*�S�VS�O]�"6�k�66����	O9܇����"����M�2J�htD1 L�\�N��25�Vbkl�f�3����s���e�En���+Z���9:��R��b������q�^����U�"5�b��yU���r���I��-iH�r����^D�bc)<��� ^�݊��J�nWM�32�]UŅ�)O���mO��Z	~]!8g���ʍZt֋�&w�!�nF��IʝsnN^K뾨8"�)�V��B�?\|�Tp &I�:�������ꪽ+<",�glF�H�BJ@KI1��Y5�UK
J	�JFt���1z�X��A}!b��,�汖�!$�d*X)j���l�Dh��p߯g�j���e���l
�|��sw��l�g�=}�M��*s(��w^����J�D LJC˷ O�96��5%/Y��q���1�j��-z�\[�>.�b�!p�^y��wj�֊%��Z`Cq�(�5��ν�0� =c�
��s�3�1�Ѩ��0�E��+��^�D�ۂ�<�#]�(�;��({�Q�]��Z�=���Tj��`� s9jZ# ��-)�+���8A`u��'�2�UiH�E�x�5�_�V��"����i���x�=T�P�[~` R&���=T#����S��P$8�0F�mVی 7&���� �X-�H}�A_�&2]l��Bs\W��]g(]^f61���|���D����Q�ǎj�+�0�HB���Z���`g�#��s�d> ꋐ�q��ު�8�c/$hQ;��B�MO��$E eL� �����D�Ux�P �(�lw^��
B7�|=�zF�-� Yx�rf�V(f�9�~x�4u:�TTX�6;:r��¢�����>��aF0c�B��{8[��l` NSq���~��{N�ҬK����K��`le@�7y��T#t�%�>�)��߃�����,MDָf���<CK���,
��Q�ܕQ����������6!ш�r	�6+ �U}���>�g ˦�����F+��@�]fF���#��u�����ɒ2��6���H�
@=�@