BZh91AY&SY�� z_�Px����߰����P����B;����i �A2��h�S�Se	�OTy4	�bh�S�%SA�CC� 4��$$M�4� �ѐh�� ����� h ��   �$�j�<�M��'��&�  h$?k� �@��J��x=��_���%fa�`��Q�9�e��B �`�1�pa"�,k�Z���v ��뫪���G�7�rɣ�ԫ&	�X�UD�2¨(4���M�?��~�m����He�͋~�+��C/��2'"��ge}1
��I!*S)��������&M�_��0ü�a������Kz�/}����]�$є����I����[E�>C�����a �qcb��д5z=�)����.4�Q�E��*��V�z�*�,���r1��Y��t�L���Utt��FcG/��51CP�ͤFM:Ӧ��]ʡS*�4��YIG�'%�pZ�2��-˻ ��'+mP��QC+3J�fWbYbղ�P��ʡiٙ&5�����B8Fh�U�����cco���`ЅV^�^r����]b׮2e3�K��a�IfD�H=$����PiY��t��GZ�&.65��׌+XV�X��,��$��^�f/dvY_���NWj���]�=^T�	���,��ߧϟ�����F���4��"ά����F����SE�Ba�A��@��Q8��Dx�F���)�q�|�gf9Ѕ�j�?hvɾa��"a�C`��!p�z��7?�'2�Ή�oZ��r���$ïUNޝ���b��;I��
^���a`�1j(��'�RO�~$L�\v.�'��%eJp�Uh��t�����ʫ���ۦ�[A��#Xč,R#X��d����PP5E/F��v$����4�L�i^�:��c*��c����*�eR���,�m�����@s�V;!	�N��Ρ4eUʫ��aS���`�5`f.�4��&��t@|�]mZ !N�&61�'�8����l9oY�-;� @B��m޹�������.P���t`��Hŕ��cFTM���Vm MW�E���Rp��]#Af����b��(!Y)L�x^C!Q\'&5��-F�B���IfZ��P��!���ΰ����VZ�5�����Z�#�r;γ�)I�0B}뵂6�I�d-� }�B�M���һ���vQ��*Ä֐�@�^$"�3g<7a�3�l흇�
S�"�V>1�T�a<&Tj���B��0Ʃ�#E�h��R���Qf�}��y3C��"�	`@k*H�Ӑ�ˬ���
3�nϴ�:���v�n��B��%�2b~Z�{1��$^ɒ:,�)�rE8P���