BZh91AY&SYRXUh l߀Px����߰����P��-�0�1��$�50M�L2F�y#j@dڃS�$� i� �2hh "�Ҟ��C�  d0&&�	�&L�&	����A��zz���觊i�hi� A� H��s�J�H�D	`�P$�z�H/��uL���j\�eD�p�ch�a"�,kv���-܉�%�_p�8�7;��gvQET��6H[�+��R��LBr�QI���'��N]M�w���3E�͎9�-:`������թC�p��)ˑ!(��@
�p�1��Q٪���0�i�v�S����m����{���f(����;#�1��@D��~�԰Qr�ȤQ�A �h�5N�+�beY��4��J�yLD��)�a0h!�k��(�#Йwr�n���F���)s͍0�D�XpD�el�X��E�P��:-�ue1�T�&����J^�N��R��t�d�(j�%ʾR�HA5aAQbu!,2bXʦ��F�r���³~x�}?H�A ��m��0B�	�aO���{8,�V���Y�"ָ�P��Ϣf����JF-�(6ϣS.sHK���px�<k���e'R����P�1KY�����Fi��[��c�l����G/S������}��%/�h�^��e�<��QH
��Ӈ��� ���*�^�m��� 񤠡�<����S1��,9����`�9u�![!� _�3 ��x������b�%'j��!�ʭ�DQ�;"�7�]��2E���Mԗ�iL�*9�%�z��T��W~&s�n��i�g��S�L׻fOѪ�P�o3�P0�X��uZJ���;[)5T���J;ƃ�2�T��S�/��yz�pAx�W��TI7�\R�U��Đ+J��<��ˌȊa�2`�
RNng���F�mR�p@m��{b��¶��.�qf(1�ø��1[����~l�KYp�)#���<�z��pxTD���U�t���Nf )��m�^3B0{����0�=��Ed4I)Q;F��y#aIܜ� @��v5�"�e�JS�g���#@�T�",�S�d ���t���P��ŀO��3yRj@�l&A�N�CL(� z��c@u����*� �f�z3n�l7+Fr�6���Liz'Ԅr���A|�9sK�4&7������ubT<T/�0�p��h! ;<����e��W �m��&���(h+�v����@d(��[����
��g�20�T��
U�re��К�-i� ��xL��I�i%�qT��a`v��A����)�\�o�r�< T�#�j�f#���䋙2Fj]����.�p� ����