BZh91AY&SY�)Z �߀Px����߰����`���" p�I�H�i2i�����L�� dё�F��~4h�T`       挘� ���F	� ���EOe&��     mU� 4h@ @ ��&!�)�e<P��z����jz�`@�vR D7� $��A �
>'���_/��Yv�,P���)/���f6���,��8�?��Z ��*�.K>@QӔ�q;ʇV����$Ei0�K"d���f��I3Z@��Py�ӝ�kj�����q��c�1�A�:��ַz��)E�D���@h����2`����/I쳤ۭ]��m��gR)`���Ĵt֥ø�2d8DH!�;;<��>UF=�j{����(;�i������7F�6�f^u��M�LЦJF.tv�Y6/(�	 T�Zw\�$��D����e�D I�$M��W���j4�0�d��6h%'�����Z�DTaW;�;������Ki��]��E�H�25]�b;>�q�`6S0̙�v�[�.���2 c�*F�(9�ƈ�4q�4B��kS!�N��Q���#�f޴���(e��Kq�}����qM.cM��Nj�Y��-k!�8S5��|0�k%-$���U��0Z"u+����kB`܉e�&�QO6lÝ2Y7�ѢBk{&�h3���[	L�(�V���Ca�jE�RѧJ��(�Owpj2�&���W���uS�7!�Ld��z^/ �31�����`�!Aۿ�O�%/���j�R�jv�]���7���6�R��#%�@�������'T3��L^�3����,X]0���M��` �B2fL���w�h��Fy��a���bu�T��ی����K���D���=o6Ŀu��`��0����(���q�ސ��R��z`<hPP��{�þ&�\ň�,9��x��>D.�`-���B�zx	�v?���v�J�>)���ܷ���AЍW[�z�Y}�[{�ݩx�fl@�����H��z�N
A�{�I�����	aEy��8���i�}���4�P�n�mg� bz�.Z�`� ��$t�eH)���f'6eF�Z���[���x��0.��1,�����Q9,���E����Z-D|!ڿ6���B�PP�8)��ޭ��(>��>�Rݑ�.�.S�g���3G�4�}*���
��P�����s�7}�7By�1�M��O���$%�.9VռNG����\�(�Qr��#
���i��6N��Є�MO���"�2�
S�g�#���EwSy�.I��l�Y���������M��|�@B���Prل�)5�E�n>�P����=չ�e{t�ȱ2F1��6�R��`��O�p#�1p�\�Z��]ђ'\��`��T'U�@m�l
�����)P�z�s��+�F2��3Ɗ�tTMbdF�j�׊�6!r���t|.,+i.�8b��[!M�4-z����O��0$.��E�&�=�5��P������m%�EL�d����DW�dv"���l{1�cޑk&H�������w$S�	B��