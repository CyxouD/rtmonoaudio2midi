BZh91AY&SYSw�S �߀Px����߰����P�:��	�QU(I!4��M�7��4S�Q��j��"��@� 4d�@ �D�� ���  ��0L@0	�h�h`ba"Bh&MOڣj4� 4&F	��IO�:I(�����H�M�����/���U6Z��E�$�0�*N _Y�x�1�t���cZ��-�Mw�]�%\�{���7}2�jZ�7Xր?�,`��S$2�/�8�8W]�;�r\��,k�AZԽ!%r�HB�j�7���$�$̘�Od���| �.��ږ����̜j/s4���LL�2���BJTʄ.TM*((�h��y��vn�˕�P����]�ɵ��]�Ň�-�e�m���H���Ea��.�h�v��c)��Q��2B�[8�ʬnvwL���W\�E�e�u�	8���25ŶR �2��;�� d2�0� �:^B�iV��@@e�y�M.�̧�%�"�BQ�Xk#'-��ы6�՗	D`����`��"VR҉*��H���?|^q�$�A+�$�@",1��1|A<�{T6M#]��^n�"��}��y��W	a %�P�Q&.����*�I�C.w!�HU1S�^�z�O��3����9u�+���a�����<�ۋ?篦%�κ���yFB�)�R/����Y	ٕLNc�x�G�%�w�x�TT��#��}���h�-�g=��W����}������g8����q�lD��E�!k�!��x�q���x�]z�] %OH���X�1�tv����z��cʒ�t��}��|bR�wt���U˄ǚ����*5 �mz)�����h�&I�p�x$Ґ4�K�a8'���z9K���� D�I����2��A���A��W�D�zɑ���U��S(���ǎ���.L�'�88��U	#TnQ���@��!�@���$տm���4���m��@}k%7e�À**��cr{�����J�%/����Md�ㅤ���u�#��/?���0�}�tEHh6fM꺪�3cE�#"i�K�	�z묐����' �l#��
�5WU�("a�Q&mu]���P#~+��Ow&%�� ��2�/�,4¬(-�2�=�==�=��ϳx�s-�#��y�C��J�c'��Ў������ـIʍ�|O�yOs3s]�jY����9�Vm�L#D�z�N�E:d�ViVt�yK���q�V�h�D���,�ꀕ��Ĕ��r�2�A��X��n����E��
��M"�C�3/ڀ��&[��l�c�G�IȻ!�;��	V3#�\�V[�٤�9b4i�qj�����]��BAM��L