BZh91AY&SYJ�i� 2_�py����߰����`_S�n��=U�AP�I��'�j�OF�S�Q��4oTmC544=M=B*�0TD�ba4� 4��i�53SFST  �      j��)�Q4��f��h5h�2sL��Lф�hшd�� A""hM���djhڣ�M��� �&��� �xnBA{(��	��B	��v� <8wJ������@2s�D�@B1"�6�Ki0��:�Wէ�@p�^%��d*�s�ǅ�:-*�y��O�Ȕy`$ [l��@  @�@6�K���.�"��kj���ӥ�>N8A#�$�0���G�dU�P )]RK��9l�h�Ga�L$30ɷٺ���8�-�K;D�h�&vH��ʂ��6S\wb�\Zh4T�L�KĦ"xxH�W�+��1II]���z.RqB�" $�j3�WS(P�MIr�&���;+6����L΀�Zf�����0D������2�.j
sX�b!�o�I�,�R�XF�K
�{(��X�b���h��=��J�p�*i-�e����٠�$�T��HK��8�^�fC2d�"
T0dE��Qbi��o�D����#=g4̐��S�<��sN�V�Y�	�h��r�Ӯ>��J��(�$Rݽ
}����f5V)p]Nd���ͮ_&�.�RM�
��1H�U��?(J%��b�@4�XUee"��1aa��W�jgS�hY���=^�}�����]z8%�m��g¿�˽��2n�'�l����l��s�#�*��7�����i �,�>.�����qAݑ�����j5����s�� 9+lv	�7pq���846$��_G�O#���[4"�_�WM�r���ork�1ؼ�*�@x�8�mK���:ڋ�㔊����ϊEIk����q�X��Q��֙�2�����{��f�@7wjg} `�a�\�%2p���N��Li-zd�tŲGY���UjD�s��n��X�i[=h4e�}5�M�1.�r��v��^+��[�G���9$��Ed��OY��,�-����j�D�D�� Z�Ŕ��=���(��3�y$V	�ꮃh$sx��Ǫ^����N������j�D�#B���v�������9�P1H:��4�Y}UJ�1��F���N D	�ﶂDPT�Jp��7U#^���*���r�g��z������`O��#R5��$�1d���M��e����C�{]�E�"R�6Jm�32�$b���{7�ic�ǩ�&K�p��4��$+�-6;�%���m��_>e�,�˂��le�7lȥB7T!�=ێjk���e�~s���侮3���2�Zk�F!y%��4;����\��7m�G6J���S��йj՞�.l1|�_y!d�H�#WJ\TV}�/�6P�AU��o)�!�N~x�� 2m�V̿�׶[:�6��2��i
?��H�
	U�5�