BZh91AY&SY�U�e �߀Px����߰����`o�����)�B�$�5=�<��G�b����zjdz��SC=Pjz JT`       jzh��4��������@ �!I�@41 ѡ�&��9�&& &#4���d�#��iO�4O�d�d�H=LA�#��!0�"�r P@�sĝ��+�$���UI�`�"�H�?�S���ch�a"�.ק�p���@��#{l">u�R�C
�o+,9&�O@(�х�t �L�eC:H���!�2O���S>���k�Ri"�4�P�:v��$2�a<�h����ܐ'MR��]q����y��I00[����kҽ��ִ�� ��io�ڪw-8Sޮz%�Ј�>��"�47�i�	j�n�/�:'Q��Z7���;���K�OFDc&�Y�t����N��l-VR���l� �EPt]5�M7]�ė��D�!X��[�t�s�N�8'
��! �h��FҮ�,�]�jC�8'%��P�a�؈+n� ��u.Q�+
]UAVXu�#!��ҫ�4�����ml)�
)��
�lɆSU!�ZfP���1�I���V��z/aRt���LeU@B��]w��u`���8Ў�r)��jB�7�����A�$�BKI$�33�E9�4u��s�mZS�z"}�t��Q�H�BD8����q�6~�4ifr�� b�aC8;�ݴBɅ��OXk� �lK'�3z���{{�O������Z�7������Q�����_���'(����)�{�@Iv}<���$���}��w�K����(񥠡��}<�O�L,ŉ$Վ�;�t��.��\446$��B�}>�<ϭ�xr\��D��S�?��\��Z�|:,̮��>�H'�K�R4��N��H� ���K��e��&s���^j;3��,w�4zm�ۚ%F�������Ь0B�hR�@�4�K��pO�I�1�ٙR�"BH�+�v��X��f��4�er��&����U5��	 �������<$G���j`�H%%�H:�ܫ��&>[I��$�܋��ټ���9�����8�̔�֩�U6($�Xba�a�{Z]�l��{�D���-�i���В7� �z�G%��F����|\���DX�����/EB\�Lh���M:���$@���m$�LR���p�U"�����)ZSPD�	UD���{
�$���`O�ә��t	 �Ȳޝ��O��t��WB������I�(f��j��h�V&H�9���N�IW���)��ќ*�I*r��}�2�Zr;�<��lK0�u�(�L#�7t�7���窗�vo�g�կƂ�ȕ�\՗�}w
��8��
��q��Y
V �9�Zt�|�ٹ�������H�5#e���t�$1IR�9��&��Pr2j:��<f�A��>�K2��Ι6vD$t��9�����]��BB�W͔