BZh91AY&SY���	 �_�Px����߰����P�8�tw�7#Lf���$SI�	��y�=4�������������3P4   � ��$�M)��oRi��#F��"����&C A��Md�2 H�14Q�LĚf����1��Q��IO� $a"C�A|"}���_�	���ɰl4	5x��7ؒ�I��k4�0�]V����@�DW���τ Y��;w�za���.P���W輻�F6;�űRS�#&�1�����]���Q[5b�p�,s��ݺ3����k���v�A�I��	%9d�H��4�o�ߪ��I�.���m����f����+=(;�4�i3�.l�!lP$�D�3Z_\�jC�+��q�) �*5Q�֦7kkW�n�o��E�9
��ڭ�c��]�u�C�C �,��[[D;�.��P�,ʏ�^�)�����8U��t٢C�!%H�AKl3"��j��$D*�0��m8*�7�����J-���LB<>�[1��s��S�E�(��"�d�|�M*Yo+#4	k�ܦ������)Cr*%!I�j�n)��W��d"ϯ���y$66����!(B��iW���/�u�^�a��R^���a5�Q�F4Ɇ�Pһ_�46*�S(b񰹾7g����i��pc�	lE��`��M'�Ru��3��q���"J�!��6��RuW?���L� pa�Ik)P%����.D�+�LEM���#�w��Ȇ�rx�o�8�ϴ�LŢ�X�ռ7��p�:�"P��́/1�3:��Pv7+�,u"4���E����9�b�J�[r�1d��%'�^L[@�)jG,R-�(���T���E���O`�,PՄ�U�ߧ`ۖy�_K����������h#�h0�Ī����{�G5�n�0���55�Z1�P���LḞÅu���W�,"��T�nRV/�J�-�hs�X��9s�L�� �D3�(�̥��,̥��K-�mÔ�d�4�3(�,u��"�B�L���u���Llc�/��q��i�ժ��s9�\0�����5�V�1�3=x�"��zAډ���t�F�0�[�i�Q8�O%nb@A5_�y�`u���3��w.���VYr�VP��)L�y^S ���N� �k��a@���a"�p��La���,������H'f�ݬ�^q�5�L��tw���%$L2�%~A�,p�!�?
���(�����੻&��U�8vJ��b 8�a��`�jN��o��+a�lMoq�Qbq�n�"����Z�	cj���pGEY!��ap��K�x�3��B�"�,H�ω{r�Ѩ���	��g���*E+�%E��q�����dQ�Ŀ�6D�jwH��$f�}����w$S�	o��