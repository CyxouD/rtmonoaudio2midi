BZh91AY&SY�B�2 G߀Px����߰����`?z�p�䦍��	$!���Sf�&ҍ�hh���ƀ���� @  �101��&%4I��4h426� �@ 44d���`F�b0L�`�!4�OM224S�l���PQ��B@����Xĉ��(HH� D	?��������m$Q@��	��H��Ą^0E�m�!�U��ut-><W�0�fd#��
X/i��R�4��>��Y(� /��@Bˮ\3�$�)CA!en�z�W]�6fq"�ՙWGj��7$���BBX�xtY��=8Z�������pٻp���k�ՠ�mL��l&׼t��dΑ䍌�]\�h�㳫��2�b������(9p8_,�m"lr(�A�Y��H D҅ݴ״,# ӄ�
R'7]��Y��|W���l
5m��cv�rh�YH�"�cS�D H�U#��[C�-E �#,Q%�,�s����pM�v���iE�`�.K0�Hg�W���ݝ`J�$!K�6��a���
E0�7Kq�@TP%�b�Z� ���	L��C�8�T���N0ڬ��)1���!*�K"��T]0z��j�zG�n\X�BBK�$�@�r'�y���o�ԕQ��4B7���V�eD����P1�jL |�&,b(���Ōӊ�
�Z�<�� f�T�MgS�ћ���Qˣ.M�2�M��^XG����w�������1YO�{o��l��S����7���ו_RFwL�򰧷���BC��Mo��2?W�i�f�4�y��5��/p��������������[�%':��!k��t��	}Z���5�;��|��ٳ�ɨ�d��[��QO��P�\�W��+f��5��r��F]Zt�(�I��;%���8�S"5ba���p s��0����z8�\JQ� 9`Y�4��+�f���3+��H�o������k����❡�h��DE8��u2�A9��6���O�K�K�����!����D�����&��9Fd�ß�d�\Uע���)����z$�@�hD�����3s�g ��i!� ��]�g��^v=�P����DUCA�A1[EBZc+"3&���hB MK�\���j�p��9��p�SUqEX�7"R%b�3��!UX��h'�Ӊ�@Ap4�S ��L���S�����C����T�0oDC٣�x�u/cH�B<�߽*Ɍe��	�p.�@>PB�]����-۞7'5/ZR�:�S��M("�X�D��O-���z��m�[�I���X�5Do��T�P0@Ἕ� �����'�Y�6B�H2�y������G��9-d%�k�K��a��l4/+�ݖ�̕U��|Fݰ9�A��<�j�b?�����秤^ɒ4��m�G���)�:	�