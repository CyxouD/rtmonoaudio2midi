BZh91AY&SY��[ |߀Px����߰����P��6�;.�5����$�L�$�4��'��ԙ<Mz��4z�T� %A h2  4d  D�BSjhi��LL@4hA��101��&$I'��Ȧ�Q���=C�SA��=A�Wl�$�X�%6"��:H�$� $�c����䭙�l�Bj�}����Q�&�ѽ�4����'"�p�[�\���h��}d<n���=Y7U�[4p��e:�;��#�;�P��p�Ȥ��K�����csh��XHeӾ�8�p�X$1�;�Ey��*a΂𛛒HJ1b��X��pk��y��j`��0��}���vr�j3��w�e�<7�	�V��g'�C[�9E��s�lr�M�63^��AVA�J��m���N��{eY����r�%�Q�QT�nP�W]�ё*�R�	r���x-3�,�Nr.�B�"�,Zl��������Q��*�i7��:��VFi��aV��+�H��{�m�uNk,3�\uKJK]5�wШ�e(�	�N,:��E¬���hg\�ԓbt�"+*EINu����ú�|����( �x��"^���w��U�#8����f�Q�Z�]1�SIP�J�ϓJ�M��+ Bb�����K�daD�ֱs�m$��X�1k_���>򓮾z�tv+��;�<~X~�_HSg�����*呶�M�iV�V�<J�Lu��W΢\r�;�@iXY��{����e��(B԰�w �G��ЋB���������m|rⰹK7�<`�ʤ��R��1�zm������K��6�;'�0H��A7+-�"DaE奝�;ĩ�-����`g��=/	2t5\c{9��vZQ��h4�U���Ht����A��b=Eg�(�ҭ�&.�O��pAx�N�X�o)Ru�MX����q�6�ե���T�`�P�p�@5��U�U�`Dn8�@�XXP-��ZF���H�c;�.���j�z﫠����a���z`�����%]=ln�t8f52@ ���8q\��ѭ��8���"�X����u��F�X&��3�uKO"jh �5=��E��-N��ԗw	�����)��E@�d�3m��!:�>��`��KѠ�\I��A�(����K�C��TX�{�m��p�kK$`:=g1�RT�!>�z�<i�86��@!:��Q��'�=g={�Z�+�$���FDdf�x�1�ҦT`�ZyEN�HY�R��TZ��hL�3U׼�+�!N�XC��,�!J���k1�pS33����H(�Ċ�e�}�&�޼kgA�>%Y���1���!Z3#�kR��Ѷ�t���#���o���"�(HGˇ-�