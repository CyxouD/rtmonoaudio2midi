BZh91AY&SYIf]m �_�Px����߰����`	�}�� B�xM�H&�����5=&T�<Bd�Oʟ�=G��L&����%@4�ɠ �@ �2b`b0#L1&L0i�	H��     hI)��?I�i�CM�z�� 4 �M=A" �1F�mG�f�FOQ�@�  4ep
���"�S0�B������9��zT��0� %�
Ƙ}e���Q ��ch��E�`��y+� Ipz���>����j5������}�z�]�]�i��щ)����E)�.i�M+�b�s��)L)�,`]RJe����N���0MI!r	�tK$v�]:m4)E�UE*�w*)�����0����ž �4E)B�o�|c��B2 �'|�%6�>��g��	�Y@2�Xm�����$�I�06?O�z4s=���w�h� ���ͺu������/G�e[%V�i���ۥxmꇔ,SRo-%�-�����2 �F�%�\�j��&�>T~_OiC�qQG��qWS�
\K�TO��퀽�훁�DjzR��ϒ@��	)�UDUj˧�f�*��X��$&FSj���w��-5�BT-ͨԑ\�V�X��T-�hc7�F�VƑ��+��2��:x��lB�9�&�i�f��[	֡zZ�Z�
EB�5t,
$����җ
���鍟"fT��dw�"�@����{.f �8�"��/�8�@���EM����q��r��������qk&b�f�e�����Q��w�1��m�>�������o{�sr����
�e���t2��AÜ�H�Y��aee��.��&&g"x	���f��V&(N�s��@������fU��T@qX�1�����)�:��p�^�([Ֆ�8݅57��\yd8���).y^_@[�
�\��WU[P�L�k����l�s�Se��U����Q����ua̮q;`�ِ��.��	�$�U.
���Lr�
�������]ܮ�eZ��O�S���g�z�oU�LŻ����|jb��Q3��w�v
���:����k����1���cH��+qd������;=�˭X�8�3*r�qSjot�:�����a"٬�:�����&v�D�����]��i�J��lÚ��3[}g5��,ty|�*�M�{����j��[���|���S���ˁ������2��͒m;G��x|�)f�JTLtH���ub�/U������\  @p  �$��m�Z��R�k�UzVyb,�g�"�Ax+tG�\\`P�Z��P��D��� �H�QPʪ�`��`eG�A�k��LeG�3�3$����ƿ��2�BQ���Wo8��>>��?O��V��L�D��yp�fڵ)$	/u�>�/�]ׂLWX�j�O�%���P<j&M�]}ǿ]�3	,��b�a���3�r$�
󔄔�y�dw�ߏk��.\}MX��;���tv��\�I����PR�Z_F=Y�C;Qdk���*.l��*0l&Z��l�s�%('n�1{�VK)o�#��C'5=�쳪�4���4��� D�`H4�\dʐS��֙#i�ɘ�ҫR�$�̧�6D�J�v�.�1L�����yYMu*T�z@�Į��6jF��l/�����0BJ�Pǆ�	�m::5��C�@��̐.F����Pl���׌زG5�\g���a�ٗ�8��G-r��͏y3D�'m� 5$	.�e���#��s�d> uE��Qz*�cE����80 S�rDPV�D���d�EwSy��$ �(�o��)`��{��`	����� IfHZ�"(;6`\(l��?��s����0A2�9�_��7�#(�r7�J/b(+8�l��҇g j	�AZn�}�:y��[3�6�&�J�쒼(a� ���J �3Zx�4�%�L�+((�Q1�Qb�m���0,^q�p`��1A[��f���z�ţ@�]t�P_���8�HxD#i�l=�~U�n��~���l�IM�'٪z3�j���"�dNc��g�u��C�V�����W/T4�ܑN$Y�[@