BZh91AY&SYW[�O �߀Px����߰����P8�q)9޴]�-j$�L�@ɪ�������'�� d=LB*�L�� LL0 �� 1B���� 4h� 4 �P�6����� &��bhb  �$
jzM��I����#L@�i���f��R�@h2
t��:�^��F-��������K�����@L!"y TSG�m���Ͳ��tC#�L���S�-Y�i�N�D�2�AI$$Zd1���?��9v0_8,���dA_��9A��Q�{�KD�p� 3��2� avՔG�<��{?Y��Ɉ�``���Ֆ^'׊���&���;�n�����sf�t<��L`�B�N�%�P��U�p�2pX0H�F�X��m4��Q��`#
Q�W(A76l�1:(���(RұCm����ˬ�н4iѻw���Wx����n��K�5Qk@���&�R�!U%��Vg���̥�%P��:Ca-tTg��e��4��("Q'�^Nlē��mTn���RM���K���ʊ�UT�8�����{�Q�a[�5%1%cD��V����{Yk��-e~y?~n!�I�O$�@""!�[����z8���|)X�Gy*�.`b0B����w��%@h�B�tD*g���恉��It�f��1`e��F�`IV�lX�=���/2r���i�3�z�y�o�	�������.�79%�!���EAb>[
 pV���G^� T<��K��G<��dG��U��~����	.������ϐ�|��ođ�)	)��X}������P���s;��Aѕ�6�c؀���愖4�����B�^��F�G!=s�0�ܱ���g;�Q)�;��I�Y<K{��'��ƒa�D=�Q�д" 5Ek �0f�Ʋ��а���27��ND'YF&.��yr��Ap���\��yQET�ˢ+�_���J(�Կ����[Y��԰w[M�lTl�ok*�GJ��ai0]�l�T?`Х1�Ġ�1kb�@}�D��͢Q���C۰���ϧÔj�F;7ؘ���r����f���+��������w��{� �n �D�2��&W���F1�[E����
�ُd�� C��P;52#1r�.���aE�j��1yLV�·�1w�Y�	�EqBK2H;��.8B�1���u����NԞ��mSV��@�{qM%'1���\m��Y��9&�x6�$��h�$u�'��̽x�+�� �1 ;=v�: �i�vB��9�W��=�R�q*J�N�,R\)Q�)	(3���HIR�IQh�&r.a��Z4
�W:CF�؎�Ǆ�pp �E�c���o�@�Φr�r(�IM���,��	%`̏y�����N�Hk�STb���@f���"�(H+����