BZh91AY&SY�<�� ,߀Px����߰����P��;!�[+VZ�I4�ړ�4�MM���bi�F!�hɠj��( �     		D���hѠ�d�4L��A�ɓ&F�L�LE�i�S�$�i��i=CF4��  �p@)�fHl$A @�RI	�M�v�Ϡ9���Vfl`�2喟�J�-ch�a�c
5ϙl��FO-���v�%�����]�n�"�?�0�ѶWL���P�2���Ŧ���x�k]V�d�ATE�b�B�WDBF1p�6[����(�$66���}�ի����~c���ʃ������l9lI���BD3"�Y^������<��`nc�z��9�
v�:������8[R�`�V�M��-A��.�8d��U�tV+*+��Z��I"�ԣ�2���82c�(,�t��S�,� Q"�dkj�%M�zj�W;��4�Qڬ������R!��i`�0�e�4^D�+��
+��^�Sbc=&vՙ#�VL3s��pq6����m��4$B���������K�Z��&L�o�{��F:cт�a~H�B�d�M��b���$1t���,�O$&L(՝e�ed� �M�M���k+�,��ve����k���c�f�?���RÿǺ����Ki�(OL��#��zv�	����ҁWuDy7����3&��oY���as1Ƅ��4��S~�� ���`��$~� m�W@����ĲQJ=*���G'�G���w��˝鄺�"Ϣ^~s�h��:�o="9����,Li��E����%z�q�%Zi2o�W8�]��n�8�m��4�IHn�J��B2y88��F�j$g�D��<�*�D�$W�Q_Ђ�W>���iU�U(/��Hп�w;H�9c���]0hH�P7c��*�*�Un_���6XKne��v�f-�h+���d}�ÒDj��E�w� $Y�;��x��Ds�Ϧ6��cD�7!,��ϩk�F�s\o{`���b&A��y$R�a�c1D�,�Eh�%�{��P� ˙�N8�7.���VXr��:*���γ��-�`CgD�=;�^����5�	���yACD'���]�ı4���'���{��^�aθ� ���"n8`���	)WmB7&E�-<!� Hr⫎�Vt��at����j�����HÊ��H�z4e��aF�R�l�t��b1����Mm�%���Y��F&	\@�6Y*"�9>���@�R��A��V���(D&i$�j=7�ܪ�w3����̚�r)�A2��@=rBEF��4+&�|�qųt ���H�Xx����H�
���