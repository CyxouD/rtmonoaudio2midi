BZh91AY&SY�76� _�Px����߰����P��6pGqF�1NH)�11�6�44�$f�=##G�<��S�i*     ������d d4� �M�	���dɓ#	�i�F& �"HѠE�OI����d Ѡ�A$�yހRa"H!%�^�w��r?����Q��l��5L>�����`���s���6���.�Vk���[c23�E��{��Ӝ�	ܺ����1�����x���B�b�_�r���<��Y`���88T�v&b���e;k�A�M��	
�� /U�~?Y��jb�0���v�}'.�s�[[M��V�_���fc*&�DtO��~5��f��gd٭i0gv=|�K��05�y8R�F�62���2ٞJ淌k)�Ԑ��1/'0٤:����EBψK��+��]Z�og2b��&.k��j	s��U ��E���EB4�G��D���cG	z<"�)���	�e�#PY�p�*XE�������h��Ŭ"�%����2J�Y&O9������7�ccoy��`�E/UN"%����N�VL���e�a����
��`�.h���>6Ķ��/ �:��½����Wѝ�L@؅{W������9QG~���+�G�����y�������|���Y�U��לfd�F�1��m���SdR��4����b#ۻ���IK��=|γ�팭�֐�6��)7��B-��G������j����ȚQ�'<~w-��;�FVp�r���"�!��^]���X��FǤF�=vd�����e�k硜�.BS�w
�'��zL�VL��>d�6.0��p��:l�5��J��� 4�C[��Td���P���b+��D�'�$̨Y�d�Pb1��~��o1q;���_��B���f�A����LB%%��J���>%>-AP�to��zI����0�Ƙ��1�dm�\�V�NX�j"4��0�Z��{g�����'��Fړ<8��.d	m�K�v��ȹ�d8��"�Q��3)���-a`����¹ŧ�64��MOf|���E�g����F�h�f�
g,�%Q��5�2�v��m}U�(�j�8�A�vR�Ct)�����!�LÓ�'����9����f���3�G#�ٵ)=�����8& ���h5��Ӌ�P���'}t�ڷF��*C�j��@�6"�3d>;Mp�3�l�G�
S�"e��t�Ob�E_¢gz��6E�O:�i��2� �uYe}��is�E�� ��T����Z��a�@�WƆr����))�l/����T3#��FLO��䋙2FʇwZ
���"�(Hm��F�