BZh91AY&SY���� O_�Px����߰����P�9.7B&�$	$��i�jbM�!��2bO!1"�       %1Dґ��Q���FM�@s F	�0M`�L$E2i&F�f)�=&��@ �F��BoI
f �H��p�x��� �_�U���`���0���"��$�"�mXCH���i^��f [%k���0�����ag�=��k�
ɚ��9,��V���a��I�L*�i�F�8�p��	��d�/�e�{�Pe
�� J�p$����U��u�0�0����G1۰5�<��5��Pp6ۚ���J9'o"Z�ᆷn�?���.sJ�
�a���d N	���ܻ�����/�}�Q�K�D�/Y����R�iLU�KC�-��f�,Q���eo��d��]��Sh��iΘp��m�@�Q���)=�����"����R{d��|�^b���B��b���2��m���ܻ�cL�F�H���Hp��3�e��7��\|���ZHHIp��HLd�ͪ�*��=��Z���H����[��Ҫ��* l�'T�EA#�ir0���nh�-\�9CsT Cd�Z�*k{]�)��OE�qY���[%���`�������8/��v�Xk𫾌O#����*@������(��b�Ǖ��6و�����F���vN�*��Ë�yn�i���?�v��Ehkhl~����&���ӭc�J=Jg���[9��:W��uze�@y�xOڗ[�l�2/zDs	�_Mt$@{,�]�������*�w��Y
��ɧ}ЄY9�vn3�d0�"Ѥ��%2k���N��L�Aަ�-\��`~3)$9�W:f{�x�V�:F2ܛi��`W�U��h�� i�
:���w�y0h2�d8%�-�7�i�)�b���9���:Iَ���Ab�/�����a�-��� (�s�k�A��#���~4K��4�+��Kps�.@,r1����XP:"�wu	�cE�F%�ԛ�P&���I`�r�����^��+:�a;�,� 2eN#J�yɄr�;O,��7E�� � -D�5��X(i�:���IR��N�=,ֹ͞�}#0p��#x�t})[,`	��Z�2\�v���9pϮP���K=����$�)(aa�$��q�B �5G^�,0�ZI0S�U8/Y`�0�2��]�J�k��𩔩���
� ��tC#E�:1d)��0�*��%׆��}�.���(�	T5���[��j로�v�ɫS�9p����T3#i�Fv%�ŝ������$h�ܖ��w$S�	���p