BZh91AY&SY� G T߀px����߰����P����'qF�,�	$�M4�MM��S��x�馡�4��cMA�~�4�   � ��0���2A�=@�4�   M �&L��L �0L�0�D����RhbI���f��  �F�!Q�ؒLH�I � h��|G�~���fd��G j0��e�+	%a�(�ѭ�4�0��yi��؀-RO������lw�xr�!��gn] �fJ�j��:���,����z�u�M�C5�v1�G�B�nk������A�)�� J��I����7�ϒI�00}��{^e�iG�~֓dX��7�wn�3�D�{�.���nQĨ��<�`�u�!��,� ����D:j(��)��`U���ܫj�=�R�{c69��ZEB�M��-P��)!@��t�c�d�U�c��.Y�Z�jSI.YdI�g����PԖ�5!��sa�Z�����J�т���� uc�q5L�)X�#��pXI�SM��15ء�s��#�8c�����R��o�͸v	 �I�IlB��IW������YZ��L2��%�C�f�TD�L軫F2&>�������@��«<y�\afaQ��]�u�����m����O�Jzi��7��?����K��_?���tc����h=*�K΋J���Hx������ ���YD	�f#ӻ���F�����1?��9�Pmv��`l������ᥡ����n��MY���{��Tw)�NZ:M�G�tg����c^H��P?�^Ll�h2t����OM����=��.�&s�?A)A;���{�
�yf�d��{��!�nc8-�2��Hm��Nw_"ӂz��j�fG���ĸ�H9g)��fX�-��4est]M�X��TS]Z�zV݂���6oL�OzpsZ�$��`����7���=+�$�VQ+�ț,k�vPZ�|4�A� Q�S����������e�cFu�\��I-���p�"���l��D����T��h��52Y6�4RDbM<�BJ	��e�P� ˙�N=��H�Y�'��YJP�D+
S9�%�0 Qg�a�Y� , ^�t��(g
��?V~������J� ���ln��`�Rd��G)�riJ�c R/���Ў�8�|2�r���1��'�]&8gU�Td�h3A'��D�A�a��cFd�+�V�S�8����S������c*,i��F��`�
U���R�#�E�Fk���{�_y �PI�MX����[y��;�g ��2k�NF�|n�
�dx(�ļ����+���&Hʷto�*��ܑN$:���