BZh91AY&SY�a�} ߀Px����߰����`>��w�9���e%p�I�*xS��	��)�hz�4�mA��E@   h   SM���24ɠ��@122i�L�)�D'�  h   ���D�����  Ѡh�H�451MLʟ�i�O�mQ�= hd]
��PB�
P����P���wF -��(��>� P�V{���ƀ��ch�a"�0kío��[1 wJ�n�X�����;��8VW3�[UI,�r�SZ�X�9QA�E
S��-�$N�qj��ҹ��ӅkA#5�ĵ�e����=r�Z�@�/m��������1 3̛���yϩl�w�[QZ�;;&��mri�4[D�`����]XP�q�
��=��se�ms �6U#�J]Ջ7�,��bvq.���Ѩ���(-#E���qhۼ:&�C1��*��K`�����>���!
.K+i��L��ˠ�$�9eT����J�H�)T��2��K�ě�m��Y�!��0৅U̫�ZUr
(,B%�^l0&�j�N>c{*ل2H�a��l�`ɉ���Q��Y^��"\����ĕw�F!)*n>��;�:�!!%}$�@� ɯB'���~����*���D�uUZ0��#�4�1�.���	g����M�Fe1Q 1rar�G~p�ax����^��`�=L���D �9�CHt��a�dS2� >��ܞg��@>CR,����,�ϳ����i� Zę�k��ו��锐ii)�a?)��D��� �z��7�9�� ѡ� $ n��'�����}D��M#��r�6��Z��N��/�ű@c� �����ia���5)����gZ�8t�{4bR߼J/N�L!$�
��*�
�;I+'4ݏ��/ql%-K��%Gp:]����A�dw���E��"D �Q]�&i���z=�4��}�D����*����%ܗgH��g_B`� �P	[U0Gev*�����G�i^VR�j���͗s(����L*b�Ƀ�R���M���s���\������'.���&vjZ@blhu��xq^ k�m~��S��@�|܋�h:9�*�S�i�I�'y5¨Ha�nU�bP�3bA	.�*e�E{���*�A5Q,��^ED�!\�� M~�K�@Oi��:D�O�\���4���NƤAC5�s]f�0mX�# �o6{R�X� �[��L�������I1Ñi��.�gU�@u�>�fzN�*�x3Rz󖾹c�
-�'�G	E�PI��Avӧ �b�^9�� ���8ۊ�2�A��Ui��1��k���B��;J$W!���4�X��]�h��j�\�՗���Q ���mW^�?OF�l�����הq��.�p�!���