BZh91AY&SY�s n߀Px����߰����P�97 �p��AXDI�1��i����4d4��A�jz �H bh ��  i��C#L�� &@  9�&& &#4���d�#��!Sl����=�=FA��=G�B %Ofa	`a" !$Ē���5�H��Y�`�Ij<�Dʈ �`�1�x0��f��Һ�{1� ]r�դ�^�-�uhUx���Hj:�g�[F�930��!��"`�Ϣ��E�cJ���,�㓅�0H�Y�)��-w_��g��	]m��B�j���]W��&����N|��������ڊ�o`�~�9�iY�<)X���I�K�k$k�@��Fl�0�D 8��F(����nq����#�b��́���ZBX��*wv`�AUh݇ԇ����F�l�J� �t@A)��!WH��b_h��I�u*�˦.WL.��)��PJ ��xC�������zS��Y4E�J��ъ�6�A�lȩ�7(ɦ�j�f�r��3$�0"n�����2H%� ��3�QN�
��٩���qނ�vDV����XL���1;�?F��VQ$	��«(;ig��	���-����
�����~�ˁ9SO�%����/w}��n�2����'����Ʃ��*�<�[0�SHm��Q��xYp!1T�c��GF��� k|�����t��*���A"�����:��`�{ ��f�/��\��y���_�b,�O4-~'L���Y��U�ˡ�Ob@�ږ�3�4LL�4A"����Ut�D�.9��&w�JqO�\�e5�/+x3���ؚ�t���pY%�ɜIĚ�9���-)�k������vԏI���Tb+)�ȷ>�͘w�ڃ1��=��S{Kc�����,
���~T".�Ƀ)��CIe�N���o�۸�ԥ�Qx-�g0�"����17 k��%��1�D�QW���{e�|��������ŚjTZ�071 t$ǵw����8��G0�#�T\CA��]EBv�1��Fe�7� �5>۳$E eKԧ �l#��
�Es���hK�d �(�}��X(U���O�#j.HD�h�AϢ���5j�<��S�=�5�~%����i�j�d�1���7�JPa�����LA�['�^�'[e�8���'~:�MQ�mK�k
��J�͡J�P���M��[�@�^�M��������T��p6wr�;7�6H� U�:s�#�Tkd)��1вׯU��p�׏9�	$ᬊF
ƾԼ�k^�'m^�Y�jŘ��IMђ�6g�A
�dvbk��1��{&H�X��?�w$S�		@ 70