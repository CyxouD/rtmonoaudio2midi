BZh91AY&SY66hF �_�Px����߰����P��ָB�V�uY����I�`����L�b�$њ����2 �H4&�(�ڞ��dɐɴM21=A��		�i�ڀbh��  ɠ��b�LFCC �#	!��?Q=OF(d�FOH F@R3��I#$Y$� PI�����ߍ����`�����Iu���bB�`���s0��F��ڻ�9��5IqF%3�v�oߤ�ukL8q>	���U����(��:�?����67liQa��j��9�Y�
�Fk�k]cǵ�`���^$"�wNK����2`�32o߉��ҵI��o��A�&�S�ۡ���ܽXv!U~�W"�:�nN�M�\V�l#&�!��Q��+V��.MU1���k�x�'2q�ggZ�V�euecEsjx2B�S���-���&�E`�t.�F*�!՜]����("�hԷ��&��hԢ(��pR��T��H'1�N�������k-0�dB��+,�z��og?'��m���Km���D!Xt�*�����u��\R`�gvK�`�d�"�|썙;08�X;�Sm+�0��ҀC���P������5�}�$������u'�8����ۗO�:��FL�e~?�wN���Յgt�g��lJ��Nu|xGG�ܣ��1<������RN��\�ƒ�����;�ϔ�L�T°r�]���������Ga���'��z��h�SqR�19u�/#�:��e��1���q��[�K���Ù�QTi�E8E%�Յ�R��O��3�P��ػ��X�a���M�*���?��_����o�)�Z$�' ;_:4��A��xK����Ґr�W�:fs-��0,��I7����*���pqO(qiDl�k���`�"RZd�K�������d;&���`[�ⴜ~!��o$-����0�g��� E2o1��D������J��fl4�R����I0�ط##�6���"ax��,!���&�h�K@�,�O�4!A5^�w
`s%I�g�#�t��Yb��2�%��������n�	��I` ���6��V(]
4H�<�=Spv�3E�l�טfK$b�擓�+f�MhF��8�a��'�W�o�/e�s�vL�Т�!���H�0Ā8vl5���F��\���00֌GR����H�Z�+�Z/*j�3��s�)�#����aa̪���1���E�� ��&�\�Y<�*�Ep���6��/V�W܋"[k���m󪯋2��l��64�;�ݬ�_�w$S�	cf�`