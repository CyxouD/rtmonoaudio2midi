BZh91AY&SY�ܳ� T_�Px����߰����P��7 �qKFL�$	$)��Oڞ����I=L�O�Fi�i�h5O�$��@    B")@�?T � 4�ѓ �`A��2`�D�M��cQ���6���h hąO,@J�  �@L^�w��8�� ���f�e ��8��[�ZI*�kF��&��5-�l�� �$���)��@�;��ZQ�a�l�l�f Ci.ڒ�[���uw������x�次��~�*�	��1r�X�ڃ������I$����9���wi�4lrv��ŏ��sς��V&ϭ]�ߋ'G>�Bo��L� HF�|��!i�XKn���@�A8t�� ���o)�t����8�GD��B-�P�Ek��DTUL�"�FH�%�iaX(f�SGb��K �(Qf�јuH��fI��a�(�r����T��"8��tv�f�s��b#s��A�WQu�l
X� �U=��v֩�!��ɭ��i��aQ('S*�jt�,������<�	�9$�@"V|E^b��z�Z^+�&YL�Ld�H>6n4�6`A���b0��V�2�9a8� ���Za�"�½����y�F�*��+k�;���Iʚ}�m�{�Go�ϖ=�ʾ����ǖ4ȴ��tȯ�F�4�+>�^EWD@����h�G�x����<h�T����a���3��������R.f������u��lo�r�Z�E	G�9���[�q�<�FW~����c�an���$���v�F�s'I��SKEB۬AcnP�^�*�:�Į�F�)IJ���z(g���mD<�oy�7(�д���UGd9�����0ZuF��&��� �b�&eyO��A��[^��o9R�ޭV.������ĎI;a��^��be�\9�J�o�F�㰇\��l��.�[�����"n��@���WKe��@(թ�a������2%~퓭�Y��,��, 8�w�u�#����\�G�h���9$R�a,�Lh�t��V�I(&�צ�B,`�Rp���F�V�s
��)�T��L���')*�z�	�p��Pbn�RA�-E��P�8�����A�ڕ
*/s���~c0l[�#��yMg��*I� �����$�Z���ؠ�Ee	�d�����m�*��3WXb 8s�z�# t�û#]�6
��g�
S�b��Js�Z��w�BE�6�@+�[�$ɷ��hɐ�BGaj�,�^�/��uĂ�9.r	V6��[�5B��K8VbQb����/6�pr��X̎�1?X���s��1d�V;���.�p�!�g�