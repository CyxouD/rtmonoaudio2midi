BZh91AY&SY��$ �߀Px����߰����Po9n��gh�Ijz���
x��ڃCj2y!��O(��
P�I�     	OQMF$G��mC#�ɍ �h4��A�ɓ&F�L�LD�	����Jy�3Қ~��4i���zGu� ���HNH�&�<�W ��ﲛ.`�"�P��bq�LIV6�L!�U��w���Zp� p���qI�ڪ6�M�m��ٍ�<t�Q#J@v蓯�N�.(L�66��1�2P���+�f̴i�9 Њ9I ��A������ϗmɀd��sxF��'=Kե�M��l��7��L�h�.�I�.&�=�(Z�Wz��Cp��B��9���yt�nt�.p:ɀ�r�,�&3��e&��q�
43]0dAs��%�����,hh�T+���:��%RId3$Ұtgk)����V��N,�Ρb�(�I�K���լ��,��K%�Wb%u����'�Gg�jTQ_j����VMzb�ʈ�i�e���Ȕ�36�ec*���� �t҉L����CF�, 1x���Nn��^�Ʌ�S�n��������7[�.�r�%YO���ߋ$��|���6�p�9)��7�Taӂ� }9�n�� b1STe'�97�?��(񥠡�,v���,Ũβ_OHt�ߐ�9{� ����!p����}|��W}���=P�s������2��Y(m +��.>��)j*��$Sp���g��D�l�z���|Į���miJ����li��J�@7_	��l�p�sJL.%Gh�)|�'�APt��/>8�)$ 9f+ѷJf��+W4F2��)M�`W�T��� ���vu�?��v݉�@zpj) ��V������n�	���e$l�ga�-����P����_d�L�i�쫠� 
_�G=>#�lv&��j�7�Oh�H`n1Xϑ�м@������P��#�A�!�ר�.��-CLh��Țu%{BD	�{m�����U�)� �t%���j�(�PD�	UD���s* T��'��$t ��Qd���@��y�h|���W>�Ԥ�3yD>���ýji�G3��ޕ�� ;c�Ԙ{8Zt k@)}s>c�wӄ��g
����c&�^$�0o9��:��i�$� �ZD�aJ���|��B@q`����� �rSOm�B42�A�s*�h�u�l����uĂ�@v�H�#ݐ��v�5I�}"�A����S�9�.���D@̎ҵ,�C�%�f59��d��;f0��]��BBg��