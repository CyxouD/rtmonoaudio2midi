BZh91AY&SY�[� V_�Px����߰����P/9lr3�j��Ih&��?Q��yL�4�f�G�LFF�P�e2Q�6�C&@� i�S$z$�� =@=@d  h0`��`ѐ��&��D�6��$l�
~�h�41��=MT�n�$�a"	!HDR�M�o^@//֪l��`�P¡�d��Ă�*����EXZ�G�m���,���Y&/�aEN�T�+�E*�%���j��k?8I���(H�[M�*q�2D.��8	�g�pNS�0C��BDOD����mz��+S68wU�?��ֺ�3�f��� �K��hs�{;D �4�6&�#���I�������F%�L��	BP�W�eъ;F�0�k�ŝ�j�j���LB���Y��bd�R�^ٱ��#1,d��la S �QUKb8B����T�H�yW��1A*�t��"(PH�+��P���$$�$�H1�m���"b<ލՋҳ��"Q�n��\�Ԡ5	�.̔�!��CDH�%�DoAXѝ�E}n3AqJ+�\�Q�lVōv�uƎ�4UW<���|V���p���W�����s~;7NZrW��琴�]9�@[�ti���W��f1�e:���þ��L$�_�=��aۚ�@�֝�����V���^ n��5���b�j �v���s�G�t�[�.��1,����v���-d�у�&�O\�m�"�J+���wWP�`��e=􅑑�e�ϙ���z�8������ĥ"9��4�Kd_8'�
����.>�E
@� ��+��n,�1Zx �c,��I7����*��P
�ke����yh�L�=���zʡi�Jyn�&�"oe)�J� ��ÁQ�B'I1��&�j��,�k�LN@L8��ǢOi�y��P�]â����c�,�D���.�`!�M�S��0�����IαR�P^G��+�sBR��Đ����' ����H������b�a��ɴ9F�x� !�A��,�t����yb����yO�.�+plM[]�Y9͚�M0r(�G�t���JTI��/܄YΠ��sn�� P������Y�5�'�e/Z�:-S���PG.�	�#���״,;H�B�
X����-�a0H�GI�H�0
H���Π+X
�qԞ���!J�ÙUm�Ɛ�T��GF#�H$O`�n��朴� d����r�'ĨQr%�_{�t+�����#ُ3ٍnrFfL�����cWB���"�(Hm-�@�