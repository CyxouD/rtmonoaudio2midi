BZh91AY&SY{�� �_�px����߰����P���pF�Z����I&S�M&OI�I�6���j44`A�~�I#     0 �BD!��h�d4=@�4h =@8ɓ&# &L �# C �Dɡ4Қy���M���  4�H���I",$=$ 䄧H���m_������X6��>���_�	
т&����D�Q�ǅ����[�bS?J����}�6�!ܭxSr��iiL���fZ��Q:Ts�cu�V��P�g���Ӧ3Vf�_l�50�q ��t��-D�B)�pӃ�a߿$�!�<o�6mg��jK�;]��o[N/L ����)!�YTW���ɔt�Fj�`6�Y�u���N��DFy�fK�+s#	���^��IcR�(,��@ơ�A�6u2�XHVQ
md{	��]j�
�(PB=��pZR`^Z��6���R�h@�h�B�(�g�U�Q��+ ��)t5n�~�L@Q8)y%�@�)�Xe����oO��g������+m���D!Xx�ʽ%���u��\2`�f�/�(��f��e�ɔF���1F&�LΦ !����H5@��+�V0�R�,�KH�\ԱSb�v�G��h��-�wϚ�W��_,�^S�����{�{�0O:vO�c�®
3� ��tym��a���&+���ri��a�IL��6x�չ��#�5jX������v��ů�'��|{�չb ��+��凐�<GB6oݡy�n�@yK�+�%�g&A�^�&�QH���7]�Z���z-���k��Ӹj�f�p�Y
��asMNC`�~&8m�a��Q��8i�@ӽ�M�n�	��N�wO��"Q�Bx����}�(�Ww�P�o�vئ�]� E���Ak�G��������r�X����Ч��*Fr�S%��@�rc�(1�z�Qxb��s���dr�SJ�&61��;`��!:�em83.���v� ��] ag{�9޷"��{A����(X�X���0�mO�hB�j�X�"�2�J���h�ۤhJ��%�2�%�
�JgE⼆Ep�X�{��h�3�H����{�� ��щ�y�:��V����u���8T�# �k8�	W0��n�#�2.߸0� ��8�5�ݪ��bT��'��Ió�H���՝Y��	�$�UҬ��_NRMJ���(D�����E��*�A�E�H��(�@�uYr�K6�-x���i@6$O �̗��h�c~ 顜���+QRr2�f���zT̏��B,K�ۦf=�rE̙#=N��)���"�(H=��s�