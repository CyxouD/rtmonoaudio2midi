BZh91AY&SYp�? ߀Px����߰����`|�� u`��H�e6�?$�Ǖ? �jy � �M4ɠj��A5*@      �2b`b0#L1&L0挘� ���F	� �I5O � �  hd  �C�"M4A�l��6��S��� ѠΘ
���Z�R`"�ت�@��x?���*Y�T@&R��(�#�� b0E��<XCH���p��c� K�U�v���
�n=��v�.氃���l�&�.�L���`�1�)MD�Kpbe>�J �*&�AIB%���_�<��M9�"�H˭�Lq�p��	l��2��,�w�(4��9"�� F�z�-��<t�2@�00a��U��#Į��$�V���evz���JaM�<�VE��RLTT.7�Τ�"��Ƃn�s�2�V�@Ω<��a5-��6�Ճ3*�]�H ��@ѱ��z�z� }�4˚&�z��8W�!V׈������L#��T�}�65�K<ɮr�����<"$�(r�҉��t�BdF�d,�&�>���|�b���\#	Q�< ЪQ�P�`�#;�s�Cc�)��V��`Uș�s����ػ���h������Y	�]�9�L��wUU�Mƫ"NP�3����.��"|<Bf��.<�+�b��wQ,l$A�=�G��N��U�Ql��9� ֈ�7���Bs52�g9�Cd$�"G��꯼]�R��\.��V]�]d-����gcFG�
.���.���ܸcY��r5����_߇�Y,lm��l!( �l�S�J_O�uUԬ�%��+T����X9b����-�[��P5-B�b�L\�T�N��0�0�0���kkci�)�[e�w�Q�%���޳�D����Ow�����wu_TK	��k�8����RH�>��2�	1UC�Y()줆���X&��]��F9��	fY���0Q�y�mBD(.2HDI��1Y��h�-�Q�t�<~���M�G��F�mڗ�c�9k�Aj�_x5k"e�eJkP�]7�ow�.�0�0^�\G����Qߕ�Lಿ���U���KP����^f}ԁ���(h�$w ӥp�E �,�����Q��� I΂�u&g�w���H�[.��ޣ�ନ�)X���h�=�#u�vl�ጔJ�P�J���U����6�xJ[4��t�06󎋛Щ�f����NKU�5�3h�%]�lc�/��:���������Bfr,@Z@���r8GC;�<�0�#����fJ.��:�c,IJ'bo` @��}�I@R�)�3�n�F�Q\�n�("B	��g3�|ŀBP��N�+�=���̐%��%�"�^9�F4O<���)�,��̩��\C����6���:G��zvjb��iMt�5&��!��'(k����Dn��nκ�%�8޴�1����%h@o3��]FXK0N�VuP�,`,����V�%�A�&5�{.H��	[-4uQ�Tf�Sq�в�=��a��E���Q"�n�?���Pͪ˦l��ہT��M�1�.�	X̎���-��=���#L���ܙB����)��!��