BZh91AY&SYR#x� �_�Px����߰����P�9\gH)@�A	�hM��=<��6h���@چ�a�� QH 2z� 4  OQ��=A�=L� h 4�`LM&L�LM2100	�e5=CM���� ���%g�$�a"	!!�$����r] %���溫0`�"�$�0縛)����f6��!�]�w�-{�c�	w�lޥ@�:t�J�Ru�Qi#Z���''Q�2��g��`
R��$*�v��;\���fi'#T͵�A�,�2����� ZE�HmQ��|�S	&`@1��,�,�_�E��1�
�M�K�7&��~<,�	�:���IJ�Fq�ܥ�+�"*�Ip�-�qu���+��^4 "i �!m@@�Mf-�lD��߁M������u�E�;8y+:����H��b6ɴӲSz��ƙ���E��2��WK�1Ul�Ȁ\*՜2�-dL��S0]�Ju6m)���҅��$[�&������˔�(�� ��VJ���mH"��b�u��"i��@�SF4��3�M����ϯ����" 0� ��3:ui�4t(f��mL�n�
Y����K	h	r�,Y��UU�PiH8�dʑPb�4X����C�e�^ۙ ��-bֹ����U����>�z)�x.��_�}��P-��>��ϟ���QC���w��zg��	r�����-ϠBL[h�W*����p��ik�Vz�gsnp�	kZ��;ۃv���cC`%���˻��㵲�Z��%/US�CS�n�H��F�t�}5� >r���|��ce�@���#�S���(�zR� �3ܹ��;���JPN꺺���Xu��/�ޝY�� ���
�g1&�`1K8J�8��iָɦ�Sd\Q�bs�DeI�$ϴ��L�yE��Eb�x��L��
���A� %2;�n(��0�^u���d	B	�!�Ρ4n�Vq�߁����@��͑`�CAi�D�c3k��r�^Ƈ8Q�K�{�q���ϟ�dl��5��	�̒��^ Q���U��ɞ�@,p4QZsA��^���m�h���D�NS�d���������#@�TN�W�PE	��f�u�, JՂx|x{�y�@	k.��Zܴ�2��b_w�V���ގҮ�E��ss��f�6H�9��۝�(0�I�i�B0�PQ���Pd�W��c��/Ϛ����ա+��j���"�9e�1��9����a�3�&��c�[b)���er�R3�a�%�����KC+e�GX{���y�����R�-���s��)
�r[�$Up�^�\�t�4�����-�Į�JnF����	ffG#ؗ���f:��􍌙#+����rE8P�R#x�