BZh91AY&SY�~+ \_�px����߰����P��7 gqF�L� I �A�=	O�<#Q�=CL����C5<��$ 24 ��  !!	��A�44� � =@sbh0�2d��`�i���!�H�2���m	�{AC�z��@�LHY~p�&  ��	.�	Gܿ����S0��F�j0�n- �6I%h�ch��Ebk��Zz����%��3���;����x���t��_�k��(�ť��f�%����~�i��3j�ٍc���HPǰ�5;�f^_P�w@��r�$�`�V*��?�y�@&``����f�a��mj��XY�� q7�G�|�&�uQ�r�&7�<hE! ���O#XQ�6P{�8ی�p��ŋ���mW��;����A�[�9h�D<��,W�Θ���cr���2��˲$J�6 �N����F��GD"�n�L�i�I^L����<�"t�E�mP�ò7��Pn�e�j�l���2r��Cj�r!'�i�j�ތ�E곪�[F�)e�Q6N����hw=_�'�sI �I�I$0V;�5^R���xn���&L���֌�DY��f��*�Lk��-�Z��� KsX7N
�#
�15f��� 	�V�⍇��󗰜��׎{���/�3��Io����B��ǧ�환���<�N5䦀^W����e�� LWc��y�G�����.�>W=n�#i���ff6���\��W���b-�l�~���鿥ï�_�9���_�uI���7>���1�$q?rK�.�9�4�:�d���t�K"=���~�s��ħ�4����'���Y�h{���j���g%���K!�p1"�ᦕN��E��xA@�)��OŅ�"H唧5��+��t��c)o�4I7yiKq�)��gՆqh����0̘1���K�O4ӕS�� 7V������`�����`���9�.mA�(��,p�� �n������#�_��6O��33 ��ڷ��z�6�P�����T���B���^4ƊH���BY�$���V\��X\�Rp�պF��Yd��eVP��)L�y/�@��M���6<h`���e�IN����[�!����t���О��w9�g��0~kK$j�aӂU�H�.���$�Z����	�=5>���K],5n�j���W�Xb	8vXdB �5ZMP��M��s��)�VZ>1��o���$<�ʗ5H6@(�Hb9���(��'�qp�*W�l�1���:sI���ET^	~�r�`�X�A��W))��6�p|  TfG������>ǳ�����$eA�X����)���1X