BZh91AY&SY �P 5߀Px����߰����`�}}�� �����-�I&����=G�jz�����z�I���* `� 	� � ���&L�20�&�db``����&&�20F� 224��$��H���Q�i�@��6����5'�j�Q�z��� � ��rd�8�L�"���#B���b��w��xg� &���~!H���$,��G6�,�{ۗw˷>��w,߱�h~~ְ^_,���{��,*��3�}AF��L"#p�$'��%&DB�3�����v��XY˔ �W	��l�ݷ?��L������~sYf㯩[���i[�Я �=x����ݕ��e^.��w�=@����y���X�3�R¾�E�T*���{K��8a�6��*R�^�)�!|�o���k��ؙ:s*�΃��J*��[��D9�|tm}�+Bp
qI�K�2p$���ʊ@��ݱ�q�]��Q�W����KT�kX����WK�qY�1F�������܄���)T��<"�����S�J�!�Tx]$2��<8��eig0�C�a�zC�J�9 �L 9�j�1�r&*�n�kK�c ��X*ׅqˉk��#%�ͬ�+!,֨BN,��g�nf�7���l�̊����3�+���p�B�j���(Ua��C�sP�������;@ � �UJ(�Z�k,��^�潶�aC�U{��#R�%D!84�Mš�� ���i��-QHb���9�;녓�j���!�h�f��쎘��b�M��~k����~�����_��O�/˥��nT�I��ʥH�No/�5ڒI4�)�>1�j��!�E9;�d��'�\�,�I�Yh�$f_p�={S8k� �n)	)���ᚸ^�I3.C��B�'��Ȏ�����/��,�)x	$Iޗ&2P4
Y:4X􈱉��L	��U݁��D�E�y���o5��6ߪf�B�i���A���ZK@� �@H4�\I� �(,��#���u�+$I!΢�6�mȿ��u|�6e���%7�̶y+*��$��^��ڈ�����=i�I$L�C�S��m��Q�IN���rPZ�Wa0�Ƃ����b����}
������H��Llc�/��:��U"r��W<tg���HL�H��\���~��/��E1�T\��Ѹ�1URw6�4^H�Q;�HB�s<eWז�DP\�Jp���H�XTWqUx�P �(�ow^e��D*��{��[AZ0	$X$��Q"^[��CD'�D{<�6Ji����N�S��*ӘfU{ܑ�z,l6�\m*�N�&��=� ��*�Qv����	1�1�^,�ΪJ���@�1 ;7V���7��{�M6�p�ON5��Ƣ�МZڕ�*v�,fX㖷�q$���E��qْ�)��J��5���͚c �ٖo��!p 9H����UBѤ�\*\&g �M�t��F+�YP{�*��D�;-�~^��Hl�SLb����M�.�p� �(�